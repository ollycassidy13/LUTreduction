
module layer0_N7_ust_3(address, data);
input wire [4:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		5'd0: data = 2'd3;
		5'd1: data = 2'd3;
		5'd2: data = 2'd3;
		5'd3: data = 2'd2;
		5'd4: data = 2'd3;
		5'd5: data = 2'd3;
		5'd6: data = 2'd3;
		5'd7: data = 2'd1;
		5'd8: data = 2'd2;
		5'd9: data = 2'd2;
		5'd10: data = 2'd2;
		5'd11: data = 2'd0;
		5'd12: data = 2'd1;
		5'd13: data = 2'd2;
		5'd14: data = 2'd1;
		5'd15: data = 2'd0;
		5'd16: data = 2'd0;
		5'd17: data = 2'd1;
		5'd18: data = 2'd0;
		5'd19: data = 2'd0;
		5'd20: data = 2'd0;
		5'd21: data = 2'd0;
		5'd22: data = 2'd0;
		5'd23: data = 2'd0;
		5'd24: data = 2'd0;
		5'd25: data = 2'd0;
		5'd26: data = 2'd0;
		5'd27: data = 2'd0;
		5'd28: data = 2'd0;
		5'd29: data = 2'd0;
		5'd30: data = 2'd0;
		5'd31: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N7_rsh_3(address, data);
input wire [0:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		1'd0: data = 2'd0;
		1'd1: data = 2'd2;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N7_lb_3(address, data);
input wire [5:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		6'd0: data = 1'd1;
		6'd1: data = 1'd1;
		6'd2: data = 1'd1;
		6'd3: data = 1'd0;
		6'd4: data = 1'd0;
		6'd5: data = 1'd0;
		6'd6: data = 1'd0;
		6'd7: data = 1'd0;
		6'd8: data = 1'd0;
		6'd9: data = 1'd1;
		6'd10: data = 1'd1;
		6'd11: data = 1'd0;
		6'd12: data = 1'd1;
		6'd13: data = 1'd0;
		6'd14: data = 1'd1;
		6'd15: data = 1'd0;
		6'd16: data = 1'd1;
		6'd17: data = 1'd0;
		6'd18: data = 1'd1;
		6'd19: data = 1'd0;
		6'd20: data = 1'd0;
		6'd21: data = 1'd0;
		6'd22: data = 1'd0;
		6'd23: data = 1'd0;
		6'd24: data = 1'd0;
		6'd25: data = 1'd0;
		6'd26: data = 1'd0;
		6'd27: data = 1'd0;
		6'd28: data = 1'd0;
		6'd29: data = 1'd0;
		6'd30: data = 1'd0;
		6'd31: data = 1'd0;
		6'd32: data = 1'd0;
		6'd33: data = 1'd0;
		6'd34: data = 1'd0;
		6'd35: data = 1'd0;
		6'd36: data = 1'd0;
		6'd37: data = 1'd0;
		6'd38: data = 1'd0;
		6'd39: data = 1'd0;
		6'd40: data = 1'd0;
		6'd41: data = 1'd0;
		6'd42: data = 1'd0;
		6'd43: data = 1'd0;
		6'd44: data = 1'd0;
		6'd45: data = 1'd0;
		6'd46: data = 1'd0;
		6'd47: data = 1'd0;
		6'd48: data = 1'd0;
		6'd49: data = 1'd0;
		6'd50: data = 1'd0;
		6'd51: data = 1'd1;
		6'd52: data = 1'd0;
		6'd53: data = 1'd0;
		6'd54: data = 1'd0;
		6'd55: data = 1'd1;
		6'd56: data = 1'd0;
		6'd57: data = 1'd0;
		6'd58: data = 1'd0;
		6'd59: data = 1'd1;
		6'd60: data = 1'd0;
		6'd61: data = 1'd0;
		6'd62: data = 1'd0;
		6'd63: data = 1'd1;
		default: data = 1'd0;
	endcase
end
endmodule

module layer0_N7_3(address, data);
input wire [5:0] address;
output reg [2:0] data;

wire [1:0] t; layer0_N7_rsh_3 rsh_3_inst(address[5:5], t);
wire [0:0] lb; layer0_N7_lb_3 lb_3_inst(address, lb);
wire [1:0] u; layer0_N7_ust_3 ust_3_inst(address[4:0], u);

always @(*) begin
	data = {(u >> t), lb};
end
endmodule

module layer0_N7_ust_2(address, data);
input wire [7:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		8'd0: data = 3'd0;
		8'd1: data = 3'd4;
		8'd2: data = 3'd0;
		8'd3: data = 3'd4;
		8'd4: data = 3'd0;
		8'd5: data = 3'd4;
		8'd6: data = 3'd0;
		8'd7: data = 3'd4;
		8'd8: data = 3'd0;
		8'd9: data = 3'd1;
		8'd10: data = 3'd0;
		8'd11: data = 3'd3;
		8'd12: data = 3'd0;
		8'd13: data = 3'd4;
		8'd14: data = 3'd0;
		8'd15: data = 3'd4;
		8'd16: data = 3'd0;
		8'd17: data = 3'd3;
		8'd18: data = 3'd0;
		8'd19: data = 3'd3;
		8'd20: data = 3'd0;
		8'd21: data = 3'd2;
		8'd22: data = 3'd0;
		8'd23: data = 3'd2;
		8'd24: data = 3'd0;
		8'd25: data = 3'd1;
		8'd26: data = 3'd0;
		8'd27: data = 3'd1;
		8'd28: data = 3'd0;
		8'd29: data = 3'd1;
		8'd30: data = 3'd0;
		8'd31: data = 3'd2;
		8'd32: data = 3'd0;
		8'd33: data = 3'd3;
		8'd34: data = 3'd0;
		8'd35: data = 3'd2;
		8'd36: data = 3'd0;
		8'd37: data = 3'd1;
		8'd38: data = 3'd0;
		8'd39: data = 3'd0;
		8'd40: data = 3'd0;
		8'd41: data = 3'd3;
		8'd42: data = 3'd0;
		8'd43: data = 3'd3;
		8'd44: data = 3'd0;
		8'd45: data = 3'd3;
		8'd46: data = 3'd0;
		8'd47: data = 3'd3;
		8'd48: data = 3'd3;
		8'd49: data = 3'd4;
		8'd50: data = 3'd3;
		8'd51: data = 3'd4;
		8'd52: data = 3'd1;
		8'd53: data = 3'd4;
		8'd54: data = 3'd0;
		8'd55: data = 3'd4;
		8'd56: data = 3'd0;
		8'd57: data = 3'd4;
		8'd58: data = 3'd0;
		8'd59: data = 3'd4;
		8'd60: data = 3'd1;
		8'd61: data = 3'd4;
		8'd62: data = 3'd1;
		8'd63: data = 3'd3;
		8'd64: data = 3'd0;
		8'd65: data = 3'd4;
		8'd66: data = 3'd0;
		8'd67: data = 3'd3;
		8'd68: data = 3'd0;
		8'd69: data = 3'd3;
		8'd70: data = 3'd0;
		8'd71: data = 3'd2;
		8'd72: data = 3'd0;
		8'd73: data = 3'd3;
		8'd74: data = 3'd0;
		8'd75: data = 3'd2;
		8'd76: data = 3'd0;
		8'd77: data = 3'd2;
		8'd78: data = 3'd0;
		8'd79: data = 3'd2;
		8'd80: data = 3'd2;
		8'd81: data = 3'd3;
		8'd82: data = 3'd2;
		8'd83: data = 3'd3;
		8'd84: data = 3'd1;
		8'd85: data = 3'd3;
		8'd86: data = 3'd0;
		8'd87: data = 3'd3;
		8'd88: data = 3'd0;
		8'd89: data = 3'd2;
		8'd90: data = 3'd1;
		8'd91: data = 3'd2;
		8'd92: data = 3'd1;
		8'd93: data = 3'd2;
		8'd94: data = 3'd1;
		8'd95: data = 3'd1;
		8'd96: data = 3'd4;
		8'd97: data = 3'd6;
		8'd98: data = 3'd3;
		8'd99: data = 3'd5;
		8'd100: data = 3'd2;
		8'd101: data = 3'd5;
		8'd102: data = 3'd0;
		8'd103: data = 3'd5;
		8'd104: data = 3'd2;
		8'd105: data = 3'd5;
		8'd106: data = 3'd1;
		8'd107: data = 3'd5;
		8'd108: data = 3'd0;
		8'd109: data = 3'd4;
		8'd110: data = 3'd0;
		8'd111: data = 3'd4;
		8'd112: data = 3'd2;
		8'd113: data = 3'd3;
		8'd114: data = 3'd1;
		8'd115: data = 3'd3;
		8'd116: data = 3'd1;
		8'd117: data = 3'd3;
		8'd118: data = 3'd0;
		8'd119: data = 3'd3;
		8'd120: data = 3'd0;
		8'd121: data = 3'd2;
		8'd122: data = 3'd0;
		8'd123: data = 3'd3;
		8'd124: data = 3'd0;
		8'd125: data = 3'd3;
		8'd126: data = 3'd0;
		8'd127: data = 3'd2;
		8'd128: data = 3'd0;
		8'd129: data = 3'd0;
		8'd130: data = 3'd0;
		8'd131: data = 3'd2;
		8'd132: data = 3'd0;
		8'd133: data = 3'd3;
		8'd134: data = 3'd0;
		8'd135: data = 3'd3;
		8'd136: data = 3'd0;
		8'd137: data = 3'd3;
		8'd138: data = 3'd0;
		8'd139: data = 3'd3;
		8'd140: data = 3'd0;
		8'd141: data = 3'd3;
		8'd142: data = 3'd0;
		8'd143: data = 3'd2;
		8'd144: data = 3'd0;
		8'd145: data = 3'd3;
		8'd146: data = 3'd0;
		8'd147: data = 3'd4;
		8'd148: data = 3'd0;
		8'd149: data = 3'd3;
		8'd150: data = 3'd0;
		8'd151: data = 3'd3;
		8'd152: data = 3'd0;
		8'd153: data = 3'd3;
		8'd154: data = 3'd0;
		8'd155: data = 3'd3;
		8'd156: data = 3'd0;
		8'd157: data = 3'd3;
		8'd158: data = 3'd1;
		8'd159: data = 3'd2;
		8'd160: data = 3'd1;
		8'd161: data = 3'd2;
		8'd162: data = 3'd1;
		8'd163: data = 3'd3;
		8'd164: data = 3'd0;
		8'd165: data = 3'd3;
		8'd166: data = 3'd0;
		8'd167: data = 3'd3;
		8'd168: data = 3'd0;
		8'd169: data = 3'd0;
		8'd170: data = 3'd0;
		8'd171: data = 3'd0;
		8'd172: data = 3'd0;
		8'd173: data = 3'd2;
		8'd174: data = 3'd0;
		8'd175: data = 3'd4;
		8'd176: data = 3'd0;
		8'd177: data = 3'd4;
		8'd178: data = 3'd0;
		8'd179: data = 3'd4;
		8'd180: data = 3'd0;
		8'd181: data = 3'd3;
		8'd182: data = 3'd0;
		8'd183: data = 3'd3;
		8'd184: data = 3'd0;
		8'd185: data = 3'd4;
		8'd186: data = 3'd0;
		8'd187: data = 3'd3;
		8'd188: data = 3'd0;
		8'd189: data = 3'd3;
		8'd190: data = 3'd0;
		8'd191: data = 3'd3;
		default: data = 3'd0;
	endcase
end
endmodule

module layer0_N7_idx_2(address, data);
input wire [5:0] address;
output reg [4:0] data;

always @(*) begin
	case(address)
		6'd0: data = 5'd0;
		6'd1: data = 5'd0;
		6'd2: data = 5'd0;
		6'd3: data = 5'd10;
		6'd4: data = 5'd4;
		6'd5: data = 5'd1;
		6'd6: data = 5'd0;
		6'd7: data = 5'd6;
		6'd8: data = 5'd11;
		6'd9: data = 5'd1;
		6'd10: data = 5'd0;
		6'd11: data = 5'd12;
		6'd12: data = 5'd2;
		6'd13: data = 5'd1;
		6'd14: data = 5'd6;
		6'd15: data = 5'd13;
		6'd16: data = 5'd7;
		6'd17: data = 5'd0;
		6'd18: data = 5'd14;
		6'd19: data = 5'd8;
		6'd20: data = 5'd15;
		6'd21: data = 5'd0;
		6'd22: data = 5'd7;
		6'd23: data = 5'd4;
		6'd24: data = 5'd0;
		6'd25: data = 5'd0;
		6'd26: data = 5'd0;
		6'd27: data = 5'd0;
		6'd28: data = 5'd0;
		6'd29: data = 5'd0;
		6'd30: data = 5'd0;
		6'd31: data = 5'd0;
		6'd32: data = 5'd0;
		6'd33: data = 5'd0;
		6'd34: data = 5'd0;
		6'd35: data = 5'd0;
		6'd36: data = 5'd0;
		6'd37: data = 5'd1;
		6'd38: data = 5'd3;
		6'd39: data = 5'd4;
		6'd40: data = 5'd0;
		6'd41: data = 5'd16;
		6'd42: data = 5'd5;
		6'd43: data = 5'd17;
		6'd44: data = 5'd3;
		6'd45: data = 5'd18;
		6'd46: data = 5'd19;
		6'd47: data = 5'd20;
		6'd48: data = 5'd21;
		6'd49: data = 5'd22;
		6'd50: data = 5'd2;
		6'd51: data = 5'd3;
		6'd52: data = 5'd1;
		6'd53: data = 5'd23;
		6'd54: data = 5'd2;
		6'd55: data = 5'd0;
		6'd56: data = 5'd0;
		6'd57: data = 5'd5;
		6'd58: data = 5'd9;
		6'd59: data = 5'd0;
		6'd60: data = 5'd0;
		6'd61: data = 5'd5;
		6'd62: data = 5'd9;
		6'd63: data = 5'd8;
		default: data = 5'd0;
	endcase
end
endmodule

module layer0_N7_rsh_2(address, data);
input wire [5:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		6'd0: data = 2'd3;
		6'd1: data = 2'd3;
		6'd2: data = 2'd3;
		6'd3: data = 2'd0;
		6'd4: data = 2'd1;
		6'd5: data = 2'd2;
		6'd6: data = 2'd2;
		6'd7: data = 2'd0;
		6'd8: data = 2'd0;
		6'd9: data = 2'd2;
		6'd10: data = 2'd2;
		6'd11: data = 2'd0;
		6'd12: data = 2'd0;
		6'd13: data = 2'd2;
		6'd14: data = 2'd1;
		6'd15: data = 2'd0;
		6'd16: data = 2'd0;
		6'd17: data = 2'd1;
		6'd18: data = 2'd0;
		6'd19: data = 2'd0;
		6'd20: data = 2'd0;
		6'd21: data = 2'd1;
		6'd22: data = 2'd1;
		6'd23: data = 2'd1;
		6'd24: data = 2'd3;
		6'd25: data = 2'd3;
		6'd26: data = 2'd3;
		6'd27: data = 2'd3;
		6'd28: data = 2'd3;
		6'd29: data = 2'd3;
		6'd30: data = 2'd3;
		6'd31: data = 2'd3;
		6'd32: data = 2'd3;
		6'd33: data = 2'd3;
		6'd34: data = 2'd3;
		6'd35: data = 2'd3;
		6'd36: data = 2'd3;
		6'd37: data = 2'd2;
		6'd38: data = 2'd0;
		6'd39: data = 2'd0;
		6'd40: data = 2'd3;
		6'd41: data = 2'd0;
		6'd42: data = 2'd0;
		6'd43: data = 2'd0;
		6'd44: data = 2'd1;
		6'd45: data = 2'd0;
		6'd46: data = 2'd0;
		6'd47: data = 2'd0;
		6'd48: data = 2'd0;
		6'd49: data = 2'd0;
		6'd50: data = 2'd0;
		6'd51: data = 2'd0;
		6'd52: data = 2'd0;
		6'd53: data = 2'd0;
		6'd54: data = 2'd0;
		6'd55: data = 2'd2;
		6'd56: data = 2'd0;
		6'd57: data = 2'd0;
		6'd58: data = 2'd0;
		6'd59: data = 2'd2;
		6'd60: data = 2'd0;
		6'd61: data = 2'd0;
		6'd62: data = 2'd0;
		6'd63: data = 2'd2;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N7_2(address, data);
input wire [8:0] address;
output reg [2:0] data;

wire [4:0] i; layer0_N7_idx_2 idx_2_inst(address[8:3], i);
wire [1:0] t; layer0_N7_rsh_2 rsh_2_inst(address[8:3], t);
wire [2:0] b; layer0_N7_3 layer0_N7_3_inst(address[8:3], b);
wire [2:0] u; layer0_N7_ust_2 ust_2_inst({i, address[2:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule

module layer0_N7_ust_1(address, data);
input wire [9:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		10'd0: data = 3'd0;
		10'd1: data = 3'd1;
		10'd2: data = 3'd1;
		10'd3: data = 3'd2;
		10'd4: data = 3'd2;
		10'd5: data = 3'd3;
		10'd6: data = 3'd3;
		10'd7: data = 3'd4;
		10'd8: data = 3'd0;
		10'd9: data = 3'd1;
		10'd10: data = 3'd2;
		10'd11: data = 3'd3;
		10'd12: data = 3'd4;
		10'd13: data = 3'd5;
		10'd14: data = 3'd6;
		10'd15: data = 3'd7;
		10'd16: data = 3'd0;
		10'd17: data = 3'd0;
		10'd18: data = 3'd0;
		10'd19: data = 3'd0;
		10'd20: data = 3'd1;
		10'd21: data = 3'd1;
		10'd22: data = 3'd2;
		10'd23: data = 3'd2;
		10'd24: data = 3'd0;
		10'd25: data = 3'd0;
		10'd26: data = 3'd0;
		10'd27: data = 3'd1;
		10'd28: data = 3'd1;
		10'd29: data = 3'd2;
		10'd30: data = 3'd2;
		10'd31: data = 3'd3;
		10'd32: data = 3'd0;
		10'd33: data = 3'd1;
		10'd34: data = 3'd1;
		10'd35: data = 3'd2;
		10'd36: data = 3'd2;
		10'd37: data = 3'd2;
		10'd38: data = 3'd3;
		10'd39: data = 3'd3;
		10'd40: data = 3'd0;
		10'd41: data = 3'd1;
		10'd42: data = 3'd2;
		10'd43: data = 3'd2;
		10'd44: data = 3'd3;
		10'd45: data = 3'd3;
		10'd46: data = 3'd3;
		10'd47: data = 3'd3;
		10'd48: data = 3'd0;
		10'd49: data = 3'd0;
		10'd50: data = 3'd1;
		10'd51: data = 3'd1;
		10'd52: data = 3'd1;
		10'd53: data = 3'd2;
		10'd54: data = 3'd2;
		10'd55: data = 3'd3;
		10'd56: data = 3'd1;
		10'd57: data = 3'd0;
		10'd58: data = 3'd0;
		10'd59: data = 3'd1;
		10'd60: data = 3'd1;
		10'd61: data = 3'd2;
		10'd62: data = 3'd2;
		10'd63: data = 3'd3;
		10'd64: data = 3'd0;
		10'd65: data = 3'd1;
		10'd66: data = 3'd1;
		10'd67: data = 3'd1;
		10'd68: data = 3'd1;
		10'd69: data = 3'd1;
		10'd70: data = 3'd1;
		10'd71: data = 3'd1;
		10'd72: data = 3'd0;
		10'd73: data = 3'd1;
		10'd74: data = 3'd1;
		10'd75: data = 3'd2;
		10'd76: data = 3'd2;
		10'd77: data = 3'd3;
		10'd78: data = 3'd3;
		10'd79: data = 3'd3;
		10'd80: data = 3'd0;
		10'd81: data = 3'd0;
		10'd82: data = 3'd0;
		10'd83: data = 3'd0;
		10'd84: data = 3'd0;
		10'd85: data = 3'd0;
		10'd86: data = 3'd1;
		10'd87: data = 3'd2;
		10'd88: data = 3'd0;
		10'd89: data = 3'd0;
		10'd90: data = 3'd0;
		10'd91: data = 3'd0;
		10'd92: data = 3'd0;
		10'd93: data = 3'd1;
		10'd94: data = 3'd2;
		10'd95: data = 3'd2;
		10'd96: data = 3'd0;
		10'd97: data = 3'd1;
		10'd98: data = 3'd2;
		10'd99: data = 3'd3;
		10'd100: data = 3'd3;
		10'd101: data = 3'd4;
		10'd102: data = 3'd4;
		10'd103: data = 3'd5;
		10'd104: data = 3'd0;
		10'd105: data = 3'd1;
		10'd106: data = 3'd1;
		10'd107: data = 3'd1;
		10'd108: data = 3'd2;
		10'd109: data = 3'd2;
		10'd110: data = 3'd3;
		10'd111: data = 3'd3;
		10'd112: data = 3'd0;
		10'd113: data = 3'd1;
		10'd114: data = 3'd1;
		10'd115: data = 3'd1;
		10'd116: data = 3'd2;
		10'd117: data = 3'd2;
		10'd118: data = 3'd2;
		10'd119: data = 3'd2;
		10'd120: data = 3'd1;
		10'd121: data = 3'd0;
		10'd122: data = 3'd0;
		10'd123: data = 3'd0;
		10'd124: data = 3'd0;
		10'd125: data = 3'd0;
		10'd126: data = 3'd1;
		10'd127: data = 3'd1;
		10'd128: data = 3'd1;
		10'd129: data = 3'd1;
		10'd130: data = 3'd1;
		10'd131: data = 3'd0;
		10'd132: data = 3'd1;
		10'd133: data = 3'd1;
		10'd134: data = 3'd2;
		10'd135: data = 3'd2;
		10'd136: data = 3'd1;
		10'd137: data = 3'd1;
		10'd138: data = 3'd0;
		10'd139: data = 3'd0;
		10'd140: data = 3'd1;
		10'd141: data = 3'd1;
		10'd142: data = 3'd2;
		10'd143: data = 3'd2;
		10'd144: data = 3'd0;
		10'd145: data = 3'd1;
		10'd146: data = 3'd1;
		10'd147: data = 3'd1;
		10'd148: data = 3'd1;
		10'd149: data = 3'd1;
		10'd150: data = 3'd2;
		10'd151: data = 3'd2;
		10'd152: data = 3'd1;
		10'd153: data = 3'd0;
		10'd154: data = 3'd0;
		10'd155: data = 3'd0;
		10'd156: data = 3'd1;
		10'd157: data = 3'd1;
		10'd158: data = 3'd2;
		10'd159: data = 3'd2;
		10'd160: data = 3'd0;
		10'd161: data = 3'd0;
		10'd162: data = 3'd0;
		10'd163: data = 3'd0;
		10'd164: data = 3'd0;
		10'd165: data = 3'd1;
		10'd166: data = 3'd2;
		10'd167: data = 3'd3;
		10'd168: data = 3'd1;
		10'd169: data = 3'd1;
		10'd170: data = 3'd1;
		10'd171: data = 3'd1;
		10'd172: data = 3'd0;
		10'd173: data = 3'd1;
		10'd174: data = 3'd1;
		10'd175: data = 3'd2;
		10'd176: data = 3'd0;
		10'd177: data = 3'd0;
		10'd178: data = 3'd0;
		10'd179: data = 3'd1;
		10'd180: data = 3'd1;
		10'd181: data = 3'd2;
		10'd182: data = 3'd2;
		10'd183: data = 3'd2;
		10'd184: data = 3'd1;
		10'd185: data = 3'd1;
		10'd186: data = 3'd1;
		10'd187: data = 3'd0;
		10'd188: data = 3'd0;
		10'd189: data = 3'd1;
		10'd190: data = 3'd1;
		10'd191: data = 3'd2;
		10'd192: data = 3'd0;
		10'd193: data = 3'd0;
		10'd194: data = 3'd1;
		10'd195: data = 3'd1;
		10'd196: data = 3'd2;
		10'd197: data = 3'd2;
		10'd198: data = 3'd2;
		10'd199: data = 3'd3;
		10'd200: data = 3'd0;
		10'd201: data = 3'd1;
		10'd202: data = 3'd1;
		10'd203: data = 3'd2;
		10'd204: data = 3'd2;
		10'd205: data = 3'd2;
		10'd206: data = 3'd2;
		10'd207: data = 3'd2;
		10'd208: data = 3'd0;
		10'd209: data = 3'd1;
		10'd210: data = 3'd1;
		10'd211: data = 3'd2;
		10'd212: data = 3'd2;
		10'd213: data = 3'd3;
		10'd214: data = 3'd4;
		10'd215: data = 3'd5;
		10'd216: data = 3'd0;
		10'd217: data = 3'd0;
		10'd218: data = 3'd1;
		10'd219: data = 3'd1;
		10'd220: data = 3'd1;
		10'd221: data = 3'd1;
		10'd222: data = 3'd1;
		10'd223: data = 3'd2;
		10'd224: data = 3'd0;
		10'd225: data = 3'd0;
		10'd226: data = 3'd0;
		10'd227: data = 3'd1;
		10'd228: data = 3'd1;
		10'd229: data = 3'd2;
		10'd230: data = 3'd3;
		10'd231: data = 3'd4;
		10'd232: data = 3'd0;
		10'd233: data = 3'd0;
		10'd234: data = 3'd1;
		10'd235: data = 3'd2;
		10'd236: data = 3'd2;
		10'd237: data = 3'd2;
		10'd238: data = 3'd3;
		10'd239: data = 3'd3;
		10'd240: data = 3'd1;
		10'd241: data = 3'd1;
		10'd242: data = 3'd0;
		10'd243: data = 3'd1;
		10'd244: data = 3'd1;
		10'd245: data = 3'd2;
		10'd246: data = 3'd2;
		10'd247: data = 3'd2;
		10'd248: data = 3'd1;
		10'd249: data = 3'd1;
		10'd250: data = 3'd1;
		10'd251: data = 3'd1;
		10'd252: data = 3'd0;
		10'd253: data = 3'd1;
		10'd254: data = 3'd1;
		10'd255: data = 3'd1;
		10'd256: data = 3'd0;
		10'd257: data = 3'd0;
		10'd258: data = 3'd0;
		10'd259: data = 3'd0;
		10'd260: data = 3'd1;
		10'd261: data = 3'd2;
		10'd262: data = 3'd2;
		10'd263: data = 3'd2;
		10'd264: data = 3'd0;
		10'd265: data = 3'd1;
		10'd266: data = 3'd2;
		10'd267: data = 3'd3;
		10'd268: data = 3'd4;
		10'd269: data = 3'd4;
		10'd270: data = 3'd5;
		10'd271: data = 3'd5;
		10'd272: data = 3'd0;
		10'd273: data = 3'd0;
		10'd274: data = 3'd0;
		10'd275: data = 3'd0;
		10'd276: data = 3'd1;
		10'd277: data = 3'd2;
		10'd278: data = 3'd2;
		10'd279: data = 3'd3;
		10'd280: data = 3'd1;
		10'd281: data = 3'd1;
		10'd282: data = 3'd0;
		10'd283: data = 3'd0;
		10'd284: data = 3'd1;
		10'd285: data = 3'd2;
		10'd286: data = 3'd2;
		10'd287: data = 3'd2;
		10'd288: data = 3'd0;
		10'd289: data = 3'd0;
		10'd290: data = 3'd1;
		10'd291: data = 3'd1;
		10'd292: data = 3'd2;
		10'd293: data = 3'd3;
		10'd294: data = 3'd3;
		10'd295: data = 3'd4;
		10'd296: data = 3'd0;
		10'd297: data = 3'd1;
		10'd298: data = 3'd1;
		10'd299: data = 3'd1;
		10'd300: data = 3'd1;
		10'd301: data = 3'd1;
		10'd302: data = 3'd1;
		10'd303: data = 3'd2;
		10'd304: data = 3'd1;
		10'd305: data = 3'd0;
		10'd306: data = 3'd0;
		10'd307: data = 3'd0;
		10'd308: data = 3'd0;
		10'd309: data = 3'd1;
		10'd310: data = 3'd1;
		10'd311: data = 3'd2;
		10'd312: data = 3'd2;
		10'd313: data = 3'd1;
		10'd314: data = 3'd0;
		10'd315: data = 3'd1;
		10'd316: data = 3'd1;
		10'd317: data = 3'd2;
		10'd318: data = 3'd3;
		10'd319: data = 3'd3;
		10'd320: data = 3'd2;
		10'd321: data = 3'd2;
		10'd322: data = 3'd1;
		10'd323: data = 3'd1;
		10'd324: data = 3'd1;
		10'd325: data = 3'd1;
		10'd326: data = 3'd0;
		10'd327: data = 3'd0;
		10'd328: data = 3'd1;
		10'd329: data = 3'd0;
		10'd330: data = 3'd0;
		10'd331: data = 3'd1;
		10'd332: data = 3'd2;
		10'd333: data = 3'd2;
		10'd334: data = 3'd3;
		10'd335: data = 3'd3;
		10'd336: data = 3'd2;
		10'd337: data = 3'd2;
		10'd338: data = 3'd1;
		10'd339: data = 3'd0;
		10'd340: data = 3'd0;
		10'd341: data = 3'd1;
		10'd342: data = 3'd1;
		10'd343: data = 3'd2;
		10'd344: data = 3'd0;
		10'd345: data = 3'd1;
		10'd346: data = 3'd1;
		10'd347: data = 3'd1;
		10'd348: data = 3'd1;
		10'd349: data = 3'd0;
		10'd350: data = 3'd1;
		10'd351: data = 3'd1;
		10'd352: data = 3'd1;
		10'd353: data = 3'd1;
		10'd354: data = 3'd2;
		10'd355: data = 3'd0;
		10'd356: data = 3'd0;
		10'd357: data = 3'd0;
		10'd358: data = 3'd0;
		10'd359: data = 3'd0;
		10'd360: data = 3'd0;
		10'd361: data = 3'd1;
		10'd362: data = 3'd1;
		10'd363: data = 3'd1;
		10'd364: data = 3'd1;
		10'd365: data = 3'd2;
		10'd366: data = 3'd2;
		10'd367: data = 3'd3;
		10'd368: data = 3'd1;
		10'd369: data = 3'd0;
		10'd370: data = 3'd1;
		10'd371: data = 3'd1;
		10'd372: data = 3'd1;
		10'd373: data = 3'd1;
		10'd374: data = 3'd2;
		10'd375: data = 3'd2;
		10'd376: data = 3'd0;
		10'd377: data = 3'd0;
		10'd378: data = 3'd1;
		10'd379: data = 3'd0;
		10'd380: data = 3'd1;
		10'd381: data = 3'd1;
		10'd382: data = 3'd1;
		10'd383: data = 3'd1;
		10'd384: data = 3'd1;
		10'd385: data = 3'd0;
		10'd386: data = 3'd0;
		10'd387: data = 3'd0;
		10'd388: data = 3'd0;
		10'd389: data = 3'd1;
		10'd390: data = 3'd2;
		10'd391: data = 3'd2;
		10'd392: data = 3'd0;
		10'd393: data = 3'd1;
		10'd394: data = 3'd1;
		10'd395: data = 3'd1;
		10'd396: data = 3'd1;
		10'd397: data = 3'd2;
		10'd398: data = 3'd2;
		10'd399: data = 3'd2;
		10'd400: data = 3'd0;
		10'd401: data = 3'd0;
		10'd402: data = 3'd1;
		10'd403: data = 3'd1;
		10'd404: data = 3'd2;
		10'd405: data = 3'd1;
		10'd406: data = 3'd1;
		10'd407: data = 3'd1;
		10'd408: data = 3'd0;
		10'd409: data = 3'd0;
		10'd410: data = 3'd1;
		10'd411: data = 3'd1;
		10'd412: data = 3'd1;
		10'd413: data = 3'd2;
		10'd414: data = 3'd3;
		10'd415: data = 3'd3;
		10'd416: data = 3'd2;
		10'd417: data = 3'd1;
		10'd418: data = 3'd0;
		10'd419: data = 3'd1;
		10'd420: data = 3'd2;
		10'd421: data = 3'd2;
		10'd422: data = 3'd3;
		10'd423: data = 3'd3;
		10'd424: data = 3'd0;
		10'd425: data = 3'd1;
		10'd426: data = 3'd1;
		10'd427: data = 3'd2;
		10'd428: data = 3'd3;
		10'd429: data = 3'd3;
		10'd430: data = 3'd4;
		10'd431: data = 3'd4;
		10'd432: data = 3'd0;
		10'd433: data = 3'd0;
		10'd434: data = 3'd1;
		10'd435: data = 3'd1;
		10'd436: data = 3'd1;
		10'd437: data = 3'd1;
		10'd438: data = 3'd2;
		10'd439: data = 3'd2;
		10'd440: data = 3'd0;
		10'd441: data = 3'd0;
		10'd442: data = 3'd1;
		10'd443: data = 3'd2;
		10'd444: data = 3'd2;
		10'd445: data = 3'd3;
		10'd446: data = 3'd3;
		10'd447: data = 3'd4;
		10'd448: data = 3'd0;
		10'd449: data = 3'd1;
		10'd450: data = 3'd1;
		10'd451: data = 3'd1;
		10'd452: data = 3'd2;
		10'd453: data = 3'd2;
		10'd454: data = 3'd2;
		10'd455: data = 3'd3;
		10'd456: data = 3'd0;
		10'd457: data = 3'd0;
		10'd458: data = 3'd0;
		10'd459: data = 3'd0;
		10'd460: data = 3'd1;
		10'd461: data = 3'd1;
		10'd462: data = 3'd2;
		10'd463: data = 3'd3;
		10'd464: data = 3'd0;
		10'd465: data = 3'd0;
		10'd466: data = 3'd0;
		10'd467: data = 3'd0;
		10'd468: data = 3'd1;
		10'd469: data = 3'd2;
		10'd470: data = 3'd2;
		10'd471: data = 3'd1;
		10'd472: data = 3'd2;
		10'd473: data = 3'd1;
		10'd474: data = 3'd1;
		10'd475: data = 3'd1;
		10'd476: data = 3'd0;
		10'd477: data = 3'd0;
		10'd478: data = 3'd0;
		10'd479: data = 3'd0;
		10'd480: data = 3'd2;
		10'd481: data = 3'd2;
		10'd482: data = 3'd2;
		10'd483: data = 3'd2;
		10'd484: data = 3'd1;
		10'd485: data = 3'd1;
		10'd486: data = 3'd1;
		10'd487: data = 3'd0;
		10'd488: data = 3'd1;
		10'd489: data = 3'd1;
		10'd490: data = 3'd1;
		10'd491: data = 3'd1;
		10'd492: data = 3'd1;
		10'd493: data = 3'd0;
		10'd494: data = 3'd0;
		10'd495: data = 3'd0;
		10'd496: data = 3'd0;
		10'd497: data = 3'd0;
		10'd498: data = 3'd1;
		10'd499: data = 3'd1;
		10'd500: data = 3'd1;
		10'd501: data = 3'd1;
		10'd502: data = 3'd0;
		10'd503: data = 3'd0;
		10'd504: data = 3'd0;
		10'd505: data = 3'd0;
		10'd506: data = 3'd0;
		10'd507: data = 3'd1;
		10'd508: data = 3'd2;
		10'd509: data = 3'd2;
		10'd510: data = 3'd1;
		10'd511: data = 3'd1;
		10'd512: data = 3'd0;
		10'd513: data = 3'd0;
		10'd514: data = 3'd0;
		10'd515: data = 3'd1;
		10'd516: data = 3'd2;
		10'd517: data = 3'd2;
		10'd518: data = 3'd3;
		10'd519: data = 3'd3;
		10'd520: data = 3'd0;
		10'd521: data = 3'd0;
		10'd522: data = 3'd0;
		10'd523: data = 3'd1;
		10'd524: data = 3'd1;
		10'd525: data = 3'd2;
		10'd526: data = 3'd3;
		10'd527: data = 3'd3;
		10'd528: data = 3'd0;
		10'd529: data = 3'd1;
		10'd530: data = 3'd1;
		10'd531: data = 3'd1;
		10'd532: data = 3'd1;
		10'd533: data = 3'd1;
		10'd534: data = 3'd1;
		10'd535: data = 3'd0;
		10'd536: data = 3'd0;
		10'd537: data = 3'd1;
		10'd538: data = 3'd1;
		10'd539: data = 3'd1;
		10'd540: data = 3'd2;
		10'd541: data = 3'd1;
		10'd542: data = 3'd1;
		10'd543: data = 3'd1;
		10'd544: data = 3'd0;
		10'd545: data = 3'd0;
		10'd546: data = 3'd1;
		10'd547: data = 3'd1;
		10'd548: data = 3'd2;
		10'd549: data = 3'd2;
		10'd550: data = 3'd2;
		10'd551: data = 3'd1;
		10'd552: data = 3'd0;
		10'd553: data = 3'd1;
		10'd554: data = 3'd1;
		10'd555: data = 3'd2;
		10'd556: data = 3'd0;
		10'd557: data = 3'd0;
		10'd558: data = 3'd0;
		10'd559: data = 3'd0;
		10'd560: data = 3'd0;
		10'd561: data = 3'd1;
		10'd562: data = 3'd1;
		10'd563: data = 3'd2;
		10'd564: data = 3'd2;
		10'd565: data = 3'd3;
		10'd566: data = 3'd2;
		10'd567: data = 3'd2;
		10'd568: data = 3'd0;
		10'd569: data = 3'd0;
		10'd570: data = 3'd1;
		10'd571: data = 3'd2;
		10'd572: data = 3'd2;
		10'd573: data = 3'd3;
		10'd574: data = 3'd3;
		10'd575: data = 3'd3;
		10'd576: data = 3'd1;
		10'd577: data = 3'd1;
		10'd578: data = 3'd1;
		10'd579: data = 3'd0;
		10'd580: data = 3'd0;
		10'd581: data = 3'd0;
		10'd582: data = 3'd1;
		10'd583: data = 3'd1;
		10'd584: data = 3'd0;
		10'd585: data = 3'd0;
		10'd586: data = 3'd1;
		10'd587: data = 3'd1;
		10'd588: data = 3'd1;
		10'd589: data = 3'd1;
		10'd590: data = 3'd0;
		10'd591: data = 3'd1;
		10'd592: data = 3'd1;
		10'd593: data = 3'd1;
		10'd594: data = 3'd0;
		10'd595: data = 3'd1;
		10'd596: data = 3'd1;
		10'd597: data = 3'd1;
		10'd598: data = 3'd2;
		10'd599: data = 3'd2;
		10'd600: data = 3'd1;
		10'd601: data = 3'd1;
		10'd602: data = 3'd2;
		10'd603: data = 3'd2;
		10'd604: data = 3'd0;
		10'd605: data = 3'd0;
		10'd606: data = 3'd0;
		10'd607: data = 3'd0;
		10'd608: data = 3'd0;
		10'd609: data = 3'd1;
		10'd610: data = 3'd1;
		10'd611: data = 3'd2;
		10'd612: data = 3'd2;
		10'd613: data = 3'd1;
		10'd614: data = 3'd0;
		10'd615: data = 3'd0;
		10'd616: data = 3'd1;
		10'd617: data = 3'd1;
		10'd618: data = 3'd0;
		10'd619: data = 3'd0;
		10'd620: data = 3'd0;
		10'd621: data = 3'd1;
		10'd622: data = 3'd2;
		10'd623: data = 3'd2;
		10'd624: data = 3'd0;
		10'd625: data = 3'd0;
		10'd626: data = 3'd1;
		10'd627: data = 3'd1;
		10'd628: data = 3'd0;
		10'd629: data = 3'd0;
		10'd630: data = 3'd1;
		10'd631: data = 3'd1;
		10'd632: data = 3'd0;
		10'd633: data = 3'd0;
		10'd634: data = 3'd1;
		10'd635: data = 3'd1;
		10'd636: data = 3'd2;
		10'd637: data = 3'd2;
		10'd638: data = 3'd3;
		10'd639: data = 3'd2;
		10'd640: data = 3'd1;
		10'd641: data = 3'd0;
		10'd642: data = 3'd0;
		10'd643: data = 3'd1;
		10'd644: data = 3'd2;
		10'd645: data = 3'd2;
		10'd646: data = 3'd2;
		10'd647: data = 3'd3;
		10'd648: data = 3'd0;
		10'd649: data = 3'd1;
		10'd650: data = 3'd1;
		10'd651: data = 3'd2;
		10'd652: data = 3'd3;
		10'd653: data = 3'd3;
		10'd654: data = 3'd2;
		10'd655: data = 3'd2;
		10'd656: data = 3'd1;
		10'd657: data = 3'd0;
		10'd658: data = 3'd0;
		10'd659: data = 3'd0;
		10'd660: data = 3'd1;
		10'd661: data = 3'd1;
		10'd662: data = 3'd2;
		10'd663: data = 3'd3;
		10'd664: data = 3'd0;
		10'd665: data = 3'd0;
		10'd666: data = 3'd1;
		10'd667: data = 3'd1;
		10'd668: data = 3'd2;
		10'd669: data = 3'd2;
		10'd670: data = 3'd1;
		10'd671: data = 3'd2;
		10'd672: data = 3'd1;
		10'd673: data = 3'd1;
		10'd674: data = 3'd0;
		10'd675: data = 3'd1;
		10'd676: data = 3'd1;
		10'd677: data = 3'd2;
		10'd678: data = 3'd2;
		10'd679: data = 3'd3;
		10'd680: data = 3'd1;
		10'd681: data = 3'd1;
		10'd682: data = 3'd1;
		10'd683: data = 3'd0;
		10'd684: data = 3'd1;
		10'd685: data = 3'd1;
		10'd686: data = 3'd1;
		10'd687: data = 3'd2;
		10'd688: data = 3'd0;
		10'd689: data = 3'd1;
		10'd690: data = 3'd1;
		10'd691: data = 3'd1;
		10'd692: data = 3'd2;
		10'd693: data = 3'd2;
		10'd694: data = 3'd3;
		10'd695: data = 3'd2;
		10'd696: data = 3'd0;
		10'd697: data = 3'd0;
		10'd698: data = 3'd1;
		10'd699: data = 3'd1;
		10'd700: data = 3'd2;
		10'd701: data = 3'd3;
		10'd702: data = 3'd3;
		10'd703: data = 3'd3;
		default: data = 3'd0;
	endcase
end
endmodule

module layer0_N7_idx_1(address, data);
input wire [8:0] address;
output reg [6:0] data;

always @(*) begin
	case(address)
		9'd0: data = 7'd0;
		9'd1: data = 7'd0;
		9'd2: data = 7'd0;
		9'd3: data = 7'd0;
		9'd4: data = 7'd0;
		9'd5: data = 7'd0;
		9'd6: data = 7'd0;
		9'd7: data = 7'd0;
		9'd8: data = 7'd0;
		9'd9: data = 7'd0;
		9'd10: data = 7'd0;
		9'd11: data = 7'd0;
		9'd12: data = 7'd0;
		9'd13: data = 7'd0;
		9'd14: data = 7'd0;
		9'd15: data = 7'd0;
		9'd16: data = 7'd0;
		9'd17: data = 7'd0;
		9'd18: data = 7'd0;
		9'd19: data = 7'd0;
		9'd20: data = 7'd0;
		9'd21: data = 7'd0;
		9'd22: data = 7'd0;
		9'd23: data = 7'd0;
		9'd24: data = 7'd0;
		9'd25: data = 7'd0;
		9'd26: data = 7'd0;
		9'd27: data = 7'd0;
		9'd28: data = 7'd3;
		9'd29: data = 7'd0;
		9'd30: data = 7'd18;
		9'd31: data = 7'd0;
		9'd32: data = 7'd0;
		9'd33: data = 7'd0;
		9'd34: data = 7'd0;
		9'd35: data = 7'd0;
		9'd36: data = 7'd0;
		9'd37: data = 7'd8;
		9'd38: data = 7'd0;
		9'd39: data = 7'd5;
		9'd40: data = 7'd0;
		9'd41: data = 7'd5;
		9'd42: data = 7'd0;
		9'd43: data = 7'd8;
		9'd44: data = 7'd0;
		9'd45: data = 7'd0;
		9'd46: data = 7'd0;
		9'd47: data = 7'd0;
		9'd48: data = 7'd0;
		9'd49: data = 7'd0;
		9'd50: data = 7'd0;
		9'd51: data = 7'd0;
		9'd52: data = 7'd0;
		9'd53: data = 7'd0;
		9'd54: data = 7'd0;
		9'd55: data = 7'd0;
		9'd56: data = 7'd2;
		9'd57: data = 7'd8;
		9'd58: data = 7'd0;
		9'd59: data = 7'd8;
		9'd60: data = 7'd45;
		9'd61: data = 7'd8;
		9'd62: data = 7'd9;
		9'd63: data = 7'd5;
		9'd64: data = 7'd46;
		9'd65: data = 7'd8;
		9'd66: data = 7'd0;
		9'd67: data = 7'd5;
		9'd68: data = 7'd0;
		9'd69: data = 7'd4;
		9'd70: data = 7'd0;
		9'd71: data = 7'd14;
		9'd72: data = 7'd0;
		9'd73: data = 7'd18;
		9'd74: data = 7'd0;
		9'd75: data = 7'd37;
		9'd76: data = 7'd0;
		9'd77: data = 7'd0;
		9'd78: data = 7'd0;
		9'd79: data = 7'd2;
		9'd80: data = 7'd0;
		9'd81: data = 7'd47;
		9'd82: data = 7'd0;
		9'd83: data = 7'd5;
		9'd84: data = 7'd0;
		9'd85: data = 7'd5;
		9'd86: data = 7'd0;
		9'd87: data = 7'd5;
		9'd88: data = 7'd2;
		9'd89: data = 7'd5;
		9'd90: data = 7'd26;
		9'd91: data = 7'd25;
		9'd92: data = 7'd3;
		9'd93: data = 7'd25;
		9'd94: data = 7'd26;
		9'd95: data = 7'd14;
		9'd96: data = 7'd19;
		9'd97: data = 7'd4;
		9'd98: data = 7'd48;
		9'd99: data = 7'd3;
		9'd100: data = 7'd38;
		9'd101: data = 7'd18;
		9'd102: data = 7'd15;
		9'd103: data = 7'd27;
		9'd104: data = 7'd0;
		9'd105: data = 7'd14;
		9'd106: data = 7'd0;
		9'd107: data = 7'd49;
		9'd108: data = 7'd0;
		9'd109: data = 7'd2;
		9'd110: data = 7'd0;
		9'd111: data = 7'd3;
		9'd112: data = 7'd0;
		9'd113: data = 7'd1;
		9'd114: data = 7'd0;
		9'd115: data = 7'd5;
		9'd116: data = 7'd37;
		9'd117: data = 7'd8;
		9'd118: data = 7'd27;
		9'd119: data = 7'd50;
		9'd120: data = 7'd12;
		9'd121: data = 7'd33;
		9'd122: data = 7'd51;
		9'd123: data = 7'd12;
		9'd124: data = 7'd28;
		9'd125: data = 7'd9;
		9'd126: data = 7'd20;
		9'd127: data = 7'd29;
		9'd128: data = 7'd39;
		9'd129: data = 7'd4;
		9'd130: data = 7'd52;
		9'd131: data = 7'd4;
		9'd132: data = 7'd19;
		9'd133: data = 7'd1;
		9'd134: data = 7'd38;
		9'd135: data = 7'd18;
		9'd136: data = 7'd15;
		9'd137: data = 7'd27;
		9'd138: data = 7'd15;
		9'd139: data = 7'd4;
		9'd140: data = 7'd15;
		9'd141: data = 7'd1;
		9'd142: data = 7'd15;
		9'd143: data = 7'd3;
		9'd144: data = 7'd0;
		9'd145: data = 7'd1;
		9'd146: data = 7'd5;
		9'd147: data = 7'd4;
		9'd148: data = 7'd4;
		9'd149: data = 7'd4;
		9'd150: data = 7'd12;
		9'd151: data = 7'd4;
		9'd152: data = 7'd1;
		9'd153: data = 7'd4;
		9'd154: data = 7'd20;
		9'd155: data = 7'd4;
		9'd156: data = 7'd10;
		9'd157: data = 7'd29;
		9'd158: data = 7'd0;
		9'd159: data = 7'd53;
		9'd160: data = 7'd19;
		9'd161: data = 7'd4;
		9'd162: data = 7'd19;
		9'd163: data = 7'd26;
		9'd164: data = 7'd30;
		9'd165: data = 7'd0;
		9'd166: data = 7'd30;
		9'd167: data = 7'd14;
		9'd168: data = 7'd16;
		9'd169: data = 7'd54;
		9'd170: data = 7'd21;
		9'd171: data = 7'd0;
		9'd172: data = 7'd31;
		9'd173: data = 7'd1;
		9'd174: data = 7'd31;
		9'd175: data = 7'd3;
		9'd176: data = 7'd39;
		9'd177: data = 7'd2;
		9'd178: data = 7'd3;
		9'd179: data = 7'd3;
		9'd180: data = 7'd2;
		9'd181: data = 7'd1;
		9'd182: data = 7'd0;
		9'd183: data = 7'd25;
		9'd184: data = 7'd0;
		9'd185: data = 7'd4;
		9'd186: data = 7'd0;
		9'd187: data = 7'd1;
		9'd188: data = 7'd0;
		9'd189: data = 7'd55;
		9'd190: data = 7'd0;
		9'd191: data = 7'd28;
		9'd192: data = 7'd0;
		9'd193: data = 7'd12;
		9'd194: data = 7'd0;
		9'd195: data = 7'd33;
		9'd196: data = 7'd0;
		9'd197: data = 7'd56;
		9'd198: data = 7'd0;
		9'd199: data = 7'd14;
		9'd200: data = 7'd0;
		9'd201: data = 7'd12;
		9'd202: data = 7'd0;
		9'd203: data = 7'd0;
		9'd204: data = 7'd0;
		9'd205: data = 7'd1;
		9'd206: data = 7'd0;
		9'd207: data = 7'd3;
		9'd208: data = 7'd0;
		9'd209: data = 7'd2;
		9'd210: data = 7'd0;
		9'd211: data = 7'd0;
		9'd212: data = 7'd0;
		9'd213: data = 7'd2;
		9'd214: data = 7'd0;
		9'd215: data = 7'd3;
		9'd216: data = 7'd0;
		9'd217: data = 7'd36;
		9'd218: data = 7'd0;
		9'd219: data = 7'd2;
		9'd220: data = 7'd0;
		9'd221: data = 7'd2;
		9'd222: data = 7'd0;
		9'd223: data = 7'd57;
		9'd224: data = 7'd0;
		9'd225: data = 7'd0;
		9'd226: data = 7'd0;
		9'd227: data = 7'd0;
		9'd228: data = 7'd0;
		9'd229: data = 7'd0;
		9'd230: data = 7'd0;
		9'd231: data = 7'd2;
		9'd232: data = 7'd0;
		9'd233: data = 7'd2;
		9'd234: data = 7'd0;
		9'd235: data = 7'd2;
		9'd236: data = 7'd0;
		9'd237: data = 7'd2;
		9'd238: data = 7'd0;
		9'd239: data = 7'd0;
		9'd240: data = 7'd0;
		9'd241: data = 7'd0;
		9'd242: data = 7'd0;
		9'd243: data = 7'd0;
		9'd244: data = 7'd0;
		9'd245: data = 7'd0;
		9'd246: data = 7'd0;
		9'd247: data = 7'd0;
		9'd248: data = 7'd0;
		9'd249: data = 7'd2;
		9'd250: data = 7'd0;
		9'd251: data = 7'd36;
		9'd252: data = 7'd0;
		9'd253: data = 7'd2;
		9'd254: data = 7'd0;
		9'd255: data = 7'd2;
		9'd256: data = 7'd0;
		9'd257: data = 7'd0;
		9'd258: data = 7'd0;
		9'd259: data = 7'd0;
		9'd260: data = 7'd0;
		9'd261: data = 7'd0;
		9'd262: data = 7'd0;
		9'd263: data = 7'd0;
		9'd264: data = 7'd0;
		9'd265: data = 7'd2;
		9'd266: data = 7'd0;
		9'd267: data = 7'd0;
		9'd268: data = 7'd0;
		9'd269: data = 7'd0;
		9'd270: data = 7'd0;
		9'd271: data = 7'd0;
		9'd272: data = 7'd0;
		9'd273: data = 7'd0;
		9'd274: data = 7'd0;
		9'd275: data = 7'd0;
		9'd276: data = 7'd0;
		9'd277: data = 7'd0;
		9'd278: data = 7'd0;
		9'd279: data = 7'd0;
		9'd280: data = 7'd0;
		9'd281: data = 7'd2;
		9'd282: data = 7'd0;
		9'd283: data = 7'd0;
		9'd284: data = 7'd0;
		9'd285: data = 7'd22;
		9'd286: data = 7'd0;
		9'd287: data = 7'd3;
		9'd288: data = 7'd0;
		9'd289: data = 7'd0;
		9'd290: data = 7'd0;
		9'd291: data = 7'd0;
		9'd292: data = 7'd0;
		9'd293: data = 7'd0;
		9'd294: data = 7'd0;
		9'd295: data = 7'd10;
		9'd296: data = 7'd0;
		9'd297: data = 7'd2;
		9'd298: data = 7'd58;
		9'd299: data = 7'd22;
		9'd300: data = 7'd32;
		9'd301: data = 7'd3;
		9'd302: data = 7'd11;
		9'd303: data = 7'd42;
		9'd304: data = 7'd11;
		9'd305: data = 7'd59;
		9'd306: data = 7'd11;
		9'd307: data = 7'd40;
		9'd308: data = 7'd10;
		9'd309: data = 7'd60;
		9'd310: data = 7'd10;
		9'd311: data = 7'd61;
		9'd312: data = 7'd10;
		9'd313: data = 7'd62;
		9'd314: data = 7'd0;
		9'd315: data = 7'd5;
		9'd316: data = 7'd0;
		9'd317: data = 7'd33;
		9'd318: data = 7'd0;
		9'd319: data = 7'd1;
		9'd320: data = 7'd0;
		9'd321: data = 7'd0;
		9'd322: data = 7'd0;
		9'd323: data = 7'd2;
		9'd324: data = 7'd0;
		9'd325: data = 7'd28;
		9'd326: data = 7'd44;
		9'd327: data = 7'd2;
		9'd328: data = 7'd63;
		9'd329: data = 7'd41;
		9'd330: data = 7'd64;
		9'd331: data = 7'd42;
		9'd332: data = 7'd65;
		9'd333: data = 7'd43;
		9'd334: data = 7'd34;
		9'd335: data = 7'd66;
		9'd336: data = 7'd34;
		9'd337: data = 7'd67;
		9'd338: data = 7'd32;
		9'd339: data = 7'd68;
		9'd340: data = 7'd32;
		9'd341: data = 7'd12;
		9'd342: data = 7'd11;
		9'd343: data = 7'd22;
		9'd344: data = 7'd11;
		9'd345: data = 7'd6;
		9'd346: data = 7'd20;
		9'd347: data = 7'd1;
		9'd348: data = 7'd10;
		9'd349: data = 7'd29;
		9'd350: data = 7'd0;
		9'd351: data = 7'd12;
		9'd352: data = 7'd40;
		9'd353: data = 7'd10;
		9'd354: data = 7'd44;
		9'd355: data = 7'd11;
		9'd356: data = 7'd69;
		9'd357: data = 7'd34;
		9'd358: data = 7'd70;
		9'd359: data = 7'd2;
		9'd360: data = 7'd71;
		9'd361: data = 7'd72;
		9'd362: data = 7'd1;
		9'd363: data = 7'd73;
		9'd364: data = 7'd1;
		9'd365: data = 7'd9;
		9'd366: data = 7'd7;
		9'd367: data = 7'd9;
		9'd368: data = 7'd7;
		9'd369: data = 7'd1;
		9'd370: data = 7'd74;
		9'd371: data = 7'd1;
		9'd372: data = 7'd17;
		9'd373: data = 7'd3;
		9'd374: data = 7'd2;
		9'd375: data = 7'd0;
		9'd376: data = 7'd2;
		9'd377: data = 7'd4;
		9'd378: data = 7'd3;
		9'd379: data = 7'd22;
		9'd380: data = 7'd35;
		9'd381: data = 7'd6;
		9'd382: data = 7'd20;
		9'd383: data = 7'd1;
		9'd384: data = 7'd75;
		9'd385: data = 7'd11;
		9'd386: data = 7'd76;
		9'd387: data = 7'd3;
		9'd388: data = 7'd9;
		9'd389: data = 7'd77;
		9'd390: data = 7'd0;
		9'd391: data = 7'd78;
		9'd392: data = 7'd1;
		9'd393: data = 7'd79;
		9'd394: data = 7'd1;
		9'd395: data = 7'd3;
		9'd396: data = 7'd80;
		9'd397: data = 7'd0;
		9'd398: data = 7'd7;
		9'd399: data = 7'd13;
		9'd400: data = 7'd30;
		9'd401: data = 7'd1;
		9'd402: data = 7'd17;
		9'd403: data = 7'd6;
		9'd404: data = 7'd16;
		9'd405: data = 7'd0;
		9'd406: data = 7'd23;
		9'd407: data = 7'd4;
		9'd408: data = 7'd0;
		9'd409: data = 7'd1;
		9'd410: data = 7'd0;
		9'd411: data = 7'd13;
		9'd412: data = 7'd2;
		9'd413: data = 7'd4;
		9'd414: data = 7'd2;
		9'd415: data = 7'd3;
		9'd416: data = 7'd81;
		9'd417: data = 7'd82;
		9'd418: data = 7'd0;
		9'd419: data = 7'd23;
		9'd420: data = 7'd0;
		9'd421: data = 7'd83;
		9'd422: data = 7'd1;
		9'd423: data = 7'd1;
		9'd424: data = 7'd1;
		9'd425: data = 7'd6;
		9'd426: data = 7'd41;
		9'd427: data = 7'd0;
		9'd428: data = 7'd7;
		9'd429: data = 7'd4;
		9'd430: data = 7'd84;
		9'd431: data = 7'd1;
		9'd432: data = 7'd17;
		9'd433: data = 7'd24;
		9'd434: data = 7'd16;
		9'd435: data = 7'd3;
		9'd436: data = 7'd85;
		9'd437: data = 7'd0;
		9'd438: data = 7'd21;
		9'd439: data = 7'd13;
		9'd440: data = 7'd0;
		9'd441: data = 7'd1;
		9'd442: data = 7'd0;
		9'd443: data = 7'd24;
		9'd444: data = 7'd0;
		9'd445: data = 7'd6;
		9'd446: data = 7'd0;
		9'd447: data = 7'd13;
		9'd448: data = 7'd0;
		9'd449: data = 7'd43;
		9'd450: data = 7'd0;
		9'd451: data = 7'd86;
		9'd452: data = 7'd87;
		9'd453: data = 7'd1;
		9'd454: data = 7'd1;
		9'd455: data = 7'd6;
		9'd456: data = 7'd1;
		9'd457: data = 7'd0;
		9'd458: data = 7'd7;
		9'd459: data = 7'd0;
		9'd460: data = 7'd7;
		9'd461: data = 7'd13;
		9'd462: data = 7'd35;
		9'd463: data = 7'd1;
		9'd464: data = 7'd17;
		9'd465: data = 7'd6;
		9'd466: data = 7'd16;
		9'd467: data = 7'd0;
		9'd468: data = 7'd23;
		9'd469: data = 7'd4;
		9'd470: data = 7'd21;
		9'd471: data = 7'd1;
		9'd472: data = 7'd0;
		9'd473: data = 7'd24;
		9'd474: data = 7'd0;
		9'd475: data = 7'd3;
		9'd476: data = 7'd0;
		9'd477: data = 7'd3;
		9'd478: data = 7'd0;
		9'd479: data = 7'd6;
		9'd480: data = 7'd0;
		9'd481: data = 7'd4;
		9'd482: data = 7'd36;
		9'd483: data = 7'd1;
		9'd484: data = 7'd1;
		9'd485: data = 7'd1;
		9'd486: data = 7'd1;
		9'd487: data = 7'd3;
		9'd488: data = 7'd7;
		9'd489: data = 7'd0;
		9'd490: data = 7'd7;
		9'd491: data = 7'd13;
		9'd492: data = 7'd35;
		9'd493: data = 7'd1;
		9'd494: data = 7'd17;
		9'd495: data = 7'd24;
		9'd496: data = 7'd16;
		9'd497: data = 7'd3;
		9'd498: data = 7'd23;
		9'd499: data = 7'd9;
		9'd500: data = 7'd21;
		9'd501: data = 7'd13;
		9'd502: data = 7'd31;
		9'd503: data = 7'd1;
		9'd504: data = 7'd0;
		9'd505: data = 7'd6;
		9'd506: data = 7'd0;
		9'd507: data = 7'd0;
		9'd508: data = 7'd0;
		9'd509: data = 7'd9;
		9'd510: data = 7'd0;
		9'd511: data = 7'd4;
		default: data = 7'd0;
	endcase
end
endmodule

module layer0_N7_rsh_1(address, data);
input wire [8:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		9'd0: data = 2'd3;
		9'd1: data = 2'd3;
		9'd2: data = 2'd3;
		9'd3: data = 2'd3;
		9'd4: data = 2'd3;
		9'd5: data = 2'd3;
		9'd6: data = 2'd3;
		9'd7: data = 2'd3;
		9'd8: data = 2'd3;
		9'd9: data = 2'd3;
		9'd10: data = 2'd3;
		9'd11: data = 2'd3;
		9'd12: data = 2'd3;
		9'd13: data = 2'd3;
		9'd14: data = 2'd3;
		9'd15: data = 2'd3;
		9'd16: data = 2'd3;
		9'd17: data = 2'd3;
		9'd18: data = 2'd3;
		9'd19: data = 2'd3;
		9'd20: data = 2'd3;
		9'd21: data = 2'd3;
		9'd22: data = 2'd3;
		9'd23: data = 2'd3;
		9'd24: data = 2'd2;
		9'd25: data = 2'd3;
		9'd26: data = 2'd2;
		9'd27: data = 2'd3;
		9'd28: data = 2'd1;
		9'd29: data = 2'd3;
		9'd30: data = 2'd0;
		9'd31: data = 2'd3;
		9'd32: data = 2'd2;
		9'd33: data = 2'd3;
		9'd34: data = 2'd3;
		9'd35: data = 2'd3;
		9'd36: data = 2'd3;
		9'd37: data = 2'd0;
		9'd38: data = 2'd3;
		9'd39: data = 2'd1;
		9'd40: data = 2'd3;
		9'd41: data = 2'd1;
		9'd42: data = 2'd3;
		9'd43: data = 2'd0;
		9'd44: data = 2'd2;
		9'd45: data = 2'd3;
		9'd46: data = 2'd3;
		9'd47: data = 2'd3;
		9'd48: data = 2'd3;
		9'd49: data = 2'd3;
		9'd50: data = 2'd3;
		9'd51: data = 2'd3;
		9'd52: data = 2'd3;
		9'd53: data = 2'd3;
		9'd54: data = 2'd3;
		9'd55: data = 2'd3;
		9'd56: data = 2'd1;
		9'd57: data = 2'd0;
		9'd58: data = 2'd2;
		9'd59: data = 2'd0;
		9'd60: data = 2'd0;
		9'd61: data = 2'd0;
		9'd62: data = 2'd0;
		9'd63: data = 2'd1;
		9'd64: data = 2'd0;
		9'd65: data = 2'd0;
		9'd66: data = 2'd2;
		9'd67: data = 2'd1;
		9'd68: data = 2'd3;
		9'd69: data = 2'd1;
		9'd70: data = 2'd3;
		9'd71: data = 2'd0;
		9'd72: data = 2'd3;
		9'd73: data = 2'd0;
		9'd74: data = 2'd3;
		9'd75: data = 2'd0;
		9'd76: data = 2'd3;
		9'd77: data = 2'd2;
		9'd78: data = 2'd3;
		9'd79: data = 2'd1;
		9'd80: data = 2'd3;
		9'd81: data = 2'd0;
		9'd82: data = 2'd3;
		9'd83: data = 2'd1;
		9'd84: data = 2'd3;
		9'd85: data = 2'd1;
		9'd86: data = 2'd3;
		9'd87: data = 2'd1;
		9'd88: data = 2'd1;
		9'd89: data = 2'd1;
		9'd90: data = 2'd1;
		9'd91: data = 2'd0;
		9'd92: data = 2'd0;
		9'd93: data = 2'd0;
		9'd94: data = 2'd0;
		9'd95: data = 2'd0;
		9'd96: data = 2'd0;
		9'd97: data = 2'd1;
		9'd98: data = 2'd0;
		9'd99: data = 2'd1;
		9'd100: data = 2'd0;
		9'd101: data = 2'd0;
		9'd102: data = 2'd0;
		9'd103: data = 2'd0;
		9'd104: data = 2'd3;
		9'd105: data = 2'd0;
		9'd106: data = 2'd3;
		9'd107: data = 2'd0;
		9'd108: data = 2'd3;
		9'd109: data = 2'd1;
		9'd110: data = 2'd3;
		9'd111: data = 2'd1;
		9'd112: data = 2'd3;
		9'd113: data = 2'd2;
		9'd114: data = 2'd3;
		9'd115: data = 2'd1;
		9'd116: data = 2'd0;
		9'd117: data = 2'd0;
		9'd118: data = 2'd0;
		9'd119: data = 2'd0;
		9'd120: data = 2'd1;
		9'd121: data = 2'd1;
		9'd122: data = 2'd0;
		9'd123: data = 2'd1;
		9'd124: data = 2'd0;
		9'd125: data = 2'd0;
		9'd126: data = 2'd0;
		9'd127: data = 2'd0;
		9'd128: data = 2'd0;
		9'd129: data = 2'd1;
		9'd130: data = 2'd0;
		9'd131: data = 2'd1;
		9'd132: data = 2'd0;
		9'd133: data = 2'd2;
		9'd134: data = 2'd0;
		9'd135: data = 2'd0;
		9'd136: data = 2'd0;
		9'd137: data = 2'd0;
		9'd138: data = 2'd0;
		9'd139: data = 2'd1;
		9'd140: data = 2'd0;
		9'd141: data = 2'd2;
		9'd142: data = 2'd0;
		9'd143: data = 2'd1;
		9'd144: data = 2'd3;
		9'd145: data = 2'd2;
		9'd146: data = 2'd1;
		9'd147: data = 2'd1;
		9'd148: data = 2'd1;
		9'd149: data = 2'd1;
		9'd150: data = 2'd1;
		9'd151: data = 2'd1;
		9'd152: data = 2'd1;
		9'd153: data = 2'd1;
		9'd154: data = 2'd0;
		9'd155: data = 2'd0;
		9'd156: data = 2'd0;
		9'd157: data = 2'd0;
		9'd158: data = 2'd2;
		9'd159: data = 2'd0;
		9'd160: data = 2'd0;
		9'd161: data = 2'd0;
		9'd162: data = 2'd0;
		9'd163: data = 2'd1;
		9'd164: data = 2'd0;
		9'd165: data = 2'd1;
		9'd166: data = 2'd0;
		9'd167: data = 2'd0;
		9'd168: data = 2'd0;
		9'd169: data = 2'd0;
		9'd170: data = 2'd0;
		9'd171: data = 2'd1;
		9'd172: data = 2'd0;
		9'd173: data = 2'd2;
		9'd174: data = 2'd0;
		9'd175: data = 2'd1;
		9'd176: data = 2'd1;
		9'd177: data = 2'd1;
		9'd178: data = 2'd1;
		9'd179: data = 2'd1;
		9'd180: data = 2'd1;
		9'd181: data = 2'd2;
		9'd182: data = 2'd2;
		9'd183: data = 2'd0;
		9'd184: data = 2'd3;
		9'd185: data = 2'd0;
		9'd186: data = 2'd3;
		9'd187: data = 2'd1;
		9'd188: data = 2'd3;
		9'd189: data = 2'd0;
		9'd190: data = 2'd3;
		9'd191: data = 2'd0;
		9'd192: data = 2'd3;
		9'd193: data = 2'd1;
		9'd194: data = 2'd3;
		9'd195: data = 2'd1;
		9'd196: data = 2'd3;
		9'd197: data = 2'd0;
		9'd198: data = 2'd3;
		9'd199: data = 2'd0;
		9'd200: data = 2'd3;
		9'd201: data = 2'd1;
		9'd202: data = 2'd3;
		9'd203: data = 2'd1;
		9'd204: data = 2'd3;
		9'd205: data = 2'd2;
		9'd206: data = 2'd3;
		9'd207: data = 2'd1;
		9'd208: data = 2'd3;
		9'd209: data = 2'd1;
		9'd210: data = 2'd3;
		9'd211: data = 2'd2;
		9'd212: data = 2'd3;
		9'd213: data = 2'd1;
		9'd214: data = 2'd3;
		9'd215: data = 2'd1;
		9'd216: data = 2'd3;
		9'd217: data = 2'd1;
		9'd218: data = 2'd3;
		9'd219: data = 2'd0;
		9'd220: data = 2'd3;
		9'd221: data = 2'd0;
		9'd222: data = 2'd3;
		9'd223: data = 2'd0;
		9'd224: data = 2'd3;
		9'd225: data = 2'd3;
		9'd226: data = 2'd3;
		9'd227: data = 2'd3;
		9'd228: data = 2'd3;
		9'd229: data = 2'd2;
		9'd230: data = 2'd3;
		9'd231: data = 2'd1;
		9'd232: data = 2'd3;
		9'd233: data = 2'd1;
		9'd234: data = 2'd3;
		9'd235: data = 2'd1;
		9'd236: data = 2'd3;
		9'd237: data = 2'd1;
		9'd238: data = 2'd3;
		9'd239: data = 2'd2;
		9'd240: data = 2'd3;
		9'd241: data = 2'd2;
		9'd242: data = 2'd3;
		9'd243: data = 2'd3;
		9'd244: data = 2'd3;
		9'd245: data = 2'd3;
		9'd246: data = 2'd3;
		9'd247: data = 2'd2;
		9'd248: data = 2'd3;
		9'd249: data = 2'd1;
		9'd250: data = 2'd3;
		9'd251: data = 2'd1;
		9'd252: data = 2'd3;
		9'd253: data = 2'd0;
		9'd254: data = 2'd3;
		9'd255: data = 2'd0;
		9'd256: data = 2'd3;
		9'd257: data = 2'd3;
		9'd258: data = 2'd3;
		9'd259: data = 2'd3;
		9'd260: data = 2'd3;
		9'd261: data = 2'd3;
		9'd262: data = 2'd3;
		9'd263: data = 2'd2;
		9'd264: data = 2'd3;
		9'd265: data = 2'd1;
		9'd266: data = 2'd3;
		9'd267: data = 2'd2;
		9'd268: data = 2'd3;
		9'd269: data = 2'd3;
		9'd270: data = 2'd3;
		9'd271: data = 2'd3;
		9'd272: data = 2'd3;
		9'd273: data = 2'd3;
		9'd274: data = 2'd3;
		9'd275: data = 2'd3;
		9'd276: data = 2'd3;
		9'd277: data = 2'd3;
		9'd278: data = 2'd3;
		9'd279: data = 2'd3;
		9'd280: data = 2'd3;
		9'd281: data = 2'd1;
		9'd282: data = 2'd3;
		9'd283: data = 2'd1;
		9'd284: data = 2'd3;
		9'd285: data = 2'd0;
		9'd286: data = 2'd3;
		9'd287: data = 2'd0;
		9'd288: data = 2'd3;
		9'd289: data = 2'd3;
		9'd290: data = 2'd3;
		9'd291: data = 2'd3;
		9'd292: data = 2'd3;
		9'd293: data = 2'd2;
		9'd294: data = 2'd3;
		9'd295: data = 2'd0;
		9'd296: data = 2'd3;
		9'd297: data = 2'd0;
		9'd298: data = 2'd0;
		9'd299: data = 2'd0;
		9'd300: data = 2'd0;
		9'd301: data = 2'd1;
		9'd302: data = 2'd0;
		9'd303: data = 2'd1;
		9'd304: data = 2'd0;
		9'd305: data = 2'd0;
		9'd306: data = 2'd0;
		9'd307: data = 2'd0;
		9'd308: data = 2'd0;
		9'd309: data = 2'd0;
		9'd310: data = 2'd0;
		9'd311: data = 2'd0;
		9'd312: data = 2'd0;
		9'd313: data = 2'd0;
		9'd314: data = 2'd2;
		9'd315: data = 2'd0;
		9'd316: data = 2'd3;
		9'd317: data = 2'd0;
		9'd318: data = 2'd3;
		9'd319: data = 2'd0;
		9'd320: data = 2'd3;
		9'd321: data = 2'd2;
		9'd322: data = 2'd3;
		9'd323: data = 2'd1;
		9'd324: data = 2'd3;
		9'd325: data = 2'd1;
		9'd326: data = 2'd1;
		9'd327: data = 2'd0;
		9'd328: data = 2'd0;
		9'd329: data = 2'd0;
		9'd330: data = 2'd0;
		9'd331: data = 2'd0;
		9'd332: data = 2'd0;
		9'd333: data = 2'd0;
		9'd334: data = 2'd0;
		9'd335: data = 2'd0;
		9'd336: data = 2'd0;
		9'd337: data = 2'd0;
		9'd338: data = 2'd0;
		9'd339: data = 2'd0;
		9'd340: data = 2'd0;
		9'd341: data = 2'd1;
		9'd342: data = 2'd0;
		9'd343: data = 2'd0;
		9'd344: data = 2'd0;
		9'd345: data = 2'd0;
		9'd346: data = 2'd0;
		9'd347: data = 2'd1;
		9'd348: data = 2'd0;
		9'd349: data = 2'd0;
		9'd350: data = 2'd2;
		9'd351: data = 2'd0;
		9'd352: data = 2'd1;
		9'd353: data = 2'd0;
		9'd354: data = 2'd0;
		9'd355: data = 2'd0;
		9'd356: data = 2'd0;
		9'd357: data = 2'd0;
		9'd358: data = 2'd0;
		9'd359: data = 2'd0;
		9'd360: data = 2'd0;
		9'd361: data = 2'd0;
		9'd362: data = 2'd1;
		9'd363: data = 2'd0;
		9'd364: data = 2'd1;
		9'd365: data = 2'd0;
		9'd366: data = 2'd0;
		9'd367: data = 2'd0;
		9'd368: data = 2'd0;
		9'd369: data = 2'd1;
		9'd370: data = 2'd0;
		9'd371: data = 2'd1;
		9'd372: data = 2'd0;
		9'd373: data = 2'd0;
		9'd374: data = 2'd1;
		9'd375: data = 2'd0;
		9'd376: data = 2'd1;
		9'd377: data = 2'd0;
		9'd378: data = 2'd1;
		9'd379: data = 2'd0;
		9'd380: data = 2'd0;
		9'd381: data = 2'd0;
		9'd382: data = 2'd0;
		9'd383: data = 2'd1;
		9'd384: data = 2'd0;
		9'd385: data = 2'd0;
		9'd386: data = 2'd0;
		9'd387: data = 2'd0;
		9'd388: data = 2'd0;
		9'd389: data = 2'd0;
		9'd390: data = 2'd0;
		9'd391: data = 2'd0;
		9'd392: data = 2'd1;
		9'd393: data = 2'd0;
		9'd394: data = 2'd1;
		9'd395: data = 2'd0;
		9'd396: data = 2'd0;
		9'd397: data = 2'd0;
		9'd398: data = 2'd0;
		9'd399: data = 2'd0;
		9'd400: data = 2'd0;
		9'd401: data = 2'd1;
		9'd402: data = 2'd0;
		9'd403: data = 2'd0;
		9'd404: data = 2'd0;
		9'd405: data = 2'd0;
		9'd406: data = 2'd0;
		9'd407: data = 2'd0;
		9'd408: data = 2'd2;
		9'd409: data = 2'd1;
		9'd410: data = 2'd2;
		9'd411: data = 2'd0;
		9'd412: data = 2'd1;
		9'd413: data = 2'd0;
		9'd414: data = 2'd1;
		9'd415: data = 2'd0;
		9'd416: data = 2'd0;
		9'd417: data = 2'd0;
		9'd418: data = 2'd0;
		9'd419: data = 2'd0;
		9'd420: data = 2'd0;
		9'd421: data = 2'd0;
		9'd422: data = 2'd1;
		9'd423: data = 2'd1;
		9'd424: data = 2'd1;
		9'd425: data = 2'd0;
		9'd426: data = 2'd0;
		9'd427: data = 2'd0;
		9'd428: data = 2'd0;
		9'd429: data = 2'd0;
		9'd430: data = 2'd0;
		9'd431: data = 2'd1;
		9'd432: data = 2'd0;
		9'd433: data = 2'd0;
		9'd434: data = 2'd0;
		9'd435: data = 2'd0;
		9'd436: data = 2'd0;
		9'd437: data = 2'd0;
		9'd438: data = 2'd0;
		9'd439: data = 2'd0;
		9'd440: data = 2'd3;
		9'd441: data = 2'd1;
		9'd442: data = 2'd3;
		9'd443: data = 2'd0;
		9'd444: data = 2'd2;
		9'd445: data = 2'd0;
		9'd446: data = 2'd2;
		9'd447: data = 2'd0;
		9'd448: data = 2'd0;
		9'd449: data = 2'd0;
		9'd450: data = 2'd0;
		9'd451: data = 2'd0;
		9'd452: data = 2'd0;
		9'd453: data = 2'd1;
		9'd454: data = 2'd1;
		9'd455: data = 2'd0;
		9'd456: data = 2'd1;
		9'd457: data = 2'd0;
		9'd458: data = 2'd0;
		9'd459: data = 2'd0;
		9'd460: data = 2'd0;
		9'd461: data = 2'd0;
		9'd462: data = 2'd0;
		9'd463: data = 2'd1;
		9'd464: data = 2'd0;
		9'd465: data = 2'd0;
		9'd466: data = 2'd0;
		9'd467: data = 2'd0;
		9'd468: data = 2'd0;
		9'd469: data = 2'd0;
		9'd470: data = 2'd0;
		9'd471: data = 2'd1;
		9'd472: data = 2'd3;
		9'd473: data = 2'd0;
		9'd474: data = 2'd3;
		9'd475: data = 2'd0;
		9'd476: data = 2'd3;
		9'd477: data = 2'd0;
		9'd478: data = 2'd3;
		9'd479: data = 2'd0;
		9'd480: data = 2'd0;
		9'd481: data = 2'd0;
		9'd482: data = 2'd0;
		9'd483: data = 2'd1;
		9'd484: data = 2'd1;
		9'd485: data = 2'd1;
		9'd486: data = 2'd1;
		9'd487: data = 2'd0;
		9'd488: data = 2'd0;
		9'd489: data = 2'd0;
		9'd490: data = 2'd0;
		9'd491: data = 2'd0;
		9'd492: data = 2'd0;
		9'd493: data = 2'd1;
		9'd494: data = 2'd0;
		9'd495: data = 2'd0;
		9'd496: data = 2'd0;
		9'd497: data = 2'd0;
		9'd498: data = 2'd0;
		9'd499: data = 2'd0;
		9'd500: data = 2'd0;
		9'd501: data = 2'd0;
		9'd502: data = 2'd0;
		9'd503: data = 2'd1;
		9'd504: data = 2'd3;
		9'd505: data = 2'd0;
		9'd506: data = 2'd3;
		9'd507: data = 2'd0;
		9'd508: data = 2'd3;
		9'd509: data = 2'd0;
		9'd510: data = 2'd3;
		9'd511: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N7_lb_1(address, data);
input wire [11:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		12'd0: data = 1'd1;
		12'd1: data = 1'd1;
		12'd2: data = 1'd1;
		12'd3: data = 1'd1;
		12'd4: data = 1'd1;
		12'd5: data = 1'd1;
		12'd6: data = 1'd1;
		12'd7: data = 1'd1;
		12'd8: data = 1'd1;
		12'd9: data = 1'd1;
		12'd10: data = 1'd1;
		12'd11: data = 1'd1;
		12'd12: data = 1'd1;
		12'd13: data = 1'd1;
		12'd14: data = 1'd1;
		12'd15: data = 1'd1;
		12'd16: data = 1'd1;
		12'd17: data = 1'd1;
		12'd18: data = 1'd1;
		12'd19: data = 1'd1;
		12'd20: data = 1'd1;
		12'd21: data = 1'd1;
		12'd22: data = 1'd1;
		12'd23: data = 1'd1;
		12'd24: data = 1'd1;
		12'd25: data = 1'd1;
		12'd26: data = 1'd1;
		12'd27: data = 1'd1;
		12'd28: data = 1'd1;
		12'd29: data = 1'd1;
		12'd30: data = 1'd1;
		12'd31: data = 1'd1;
		12'd32: data = 1'd1;
		12'd33: data = 1'd1;
		12'd34: data = 1'd1;
		12'd35: data = 1'd1;
		12'd36: data = 1'd1;
		12'd37: data = 1'd1;
		12'd38: data = 1'd1;
		12'd39: data = 1'd1;
		12'd40: data = 1'd1;
		12'd41: data = 1'd1;
		12'd42: data = 1'd1;
		12'd43: data = 1'd1;
		12'd44: data = 1'd1;
		12'd45: data = 1'd1;
		12'd46: data = 1'd1;
		12'd47: data = 1'd1;
		12'd48: data = 1'd1;
		12'd49: data = 1'd1;
		12'd50: data = 1'd1;
		12'd51: data = 1'd1;
		12'd52: data = 1'd1;
		12'd53: data = 1'd1;
		12'd54: data = 1'd1;
		12'd55: data = 1'd1;
		12'd56: data = 1'd1;
		12'd57: data = 1'd1;
		12'd58: data = 1'd1;
		12'd59: data = 1'd1;
		12'd60: data = 1'd1;
		12'd61: data = 1'd1;
		12'd62: data = 1'd1;
		12'd63: data = 1'd1;
		12'd64: data = 1'd1;
		12'd65: data = 1'd1;
		12'd66: data = 1'd1;
		12'd67: data = 1'd1;
		12'd68: data = 1'd1;
		12'd69: data = 1'd1;
		12'd70: data = 1'd1;
		12'd71: data = 1'd1;
		12'd72: data = 1'd1;
		12'd73: data = 1'd1;
		12'd74: data = 1'd1;
		12'd75: data = 1'd1;
		12'd76: data = 1'd1;
		12'd77: data = 1'd1;
		12'd78: data = 1'd1;
		12'd79: data = 1'd1;
		12'd80: data = 1'd0;
		12'd81: data = 1'd1;
		12'd82: data = 1'd1;
		12'd83: data = 1'd1;
		12'd84: data = 1'd1;
		12'd85: data = 1'd1;
		12'd86: data = 1'd1;
		12'd87: data = 1'd1;
		12'd88: data = 1'd1;
		12'd89: data = 1'd1;
		12'd90: data = 1'd1;
		12'd91: data = 1'd1;
		12'd92: data = 1'd1;
		12'd93: data = 1'd1;
		12'd94: data = 1'd1;
		12'd95: data = 1'd1;
		12'd96: data = 1'd0;
		12'd97: data = 1'd0;
		12'd98: data = 1'd1;
		12'd99: data = 1'd1;
		12'd100: data = 1'd1;
		12'd101: data = 1'd1;
		12'd102: data = 1'd1;
		12'd103: data = 1'd1;
		12'd104: data = 1'd1;
		12'd105: data = 1'd1;
		12'd106: data = 1'd1;
		12'd107: data = 1'd1;
		12'd108: data = 1'd1;
		12'd109: data = 1'd1;
		12'd110: data = 1'd1;
		12'd111: data = 1'd1;
		12'd112: data = 1'd0;
		12'd113: data = 1'd0;
		12'd114: data = 1'd1;
		12'd115: data = 1'd1;
		12'd116: data = 1'd1;
		12'd117: data = 1'd1;
		12'd118: data = 1'd1;
		12'd119: data = 1'd1;
		12'd120: data = 1'd1;
		12'd121: data = 1'd1;
		12'd122: data = 1'd1;
		12'd123: data = 1'd1;
		12'd124: data = 1'd1;
		12'd125: data = 1'd1;
		12'd126: data = 1'd1;
		12'd127: data = 1'd1;
		12'd128: data = 1'd0;
		12'd129: data = 1'd0;
		12'd130: data = 1'd0;
		12'd131: data = 1'd1;
		12'd132: data = 1'd1;
		12'd133: data = 1'd1;
		12'd134: data = 1'd1;
		12'd135: data = 1'd1;
		12'd136: data = 1'd1;
		12'd137: data = 1'd1;
		12'd138: data = 1'd1;
		12'd139: data = 1'd1;
		12'd140: data = 1'd1;
		12'd141: data = 1'd1;
		12'd142: data = 1'd1;
		12'd143: data = 1'd1;
		12'd144: data = 1'd0;
		12'd145: data = 1'd0;
		12'd146: data = 1'd0;
		12'd147: data = 1'd0;
		12'd148: data = 1'd1;
		12'd149: data = 1'd1;
		12'd150: data = 1'd1;
		12'd151: data = 1'd1;
		12'd152: data = 1'd1;
		12'd153: data = 1'd1;
		12'd154: data = 1'd1;
		12'd155: data = 1'd1;
		12'd156: data = 1'd1;
		12'd157: data = 1'd1;
		12'd158: data = 1'd1;
		12'd159: data = 1'd1;
		12'd160: data = 1'd0;
		12'd161: data = 1'd0;
		12'd162: data = 1'd0;
		12'd163: data = 1'd0;
		12'd164: data = 1'd0;
		12'd165: data = 1'd1;
		12'd166: data = 1'd1;
		12'd167: data = 1'd1;
		12'd168: data = 1'd1;
		12'd169: data = 1'd1;
		12'd170: data = 1'd1;
		12'd171: data = 1'd1;
		12'd172: data = 1'd1;
		12'd173: data = 1'd1;
		12'd174: data = 1'd1;
		12'd175: data = 1'd1;
		12'd176: data = 1'd0;
		12'd177: data = 1'd0;
		12'd178: data = 1'd0;
		12'd179: data = 1'd0;
		12'd180: data = 1'd0;
		12'd181: data = 1'd0;
		12'd182: data = 1'd0;
		12'd183: data = 1'd0;
		12'd184: data = 1'd1;
		12'd185: data = 1'd1;
		12'd186: data = 1'd1;
		12'd187: data = 1'd1;
		12'd188: data = 1'd1;
		12'd189: data = 1'd1;
		12'd190: data = 1'd1;
		12'd191: data = 1'd1;
		12'd192: data = 1'd1;
		12'd193: data = 1'd1;
		12'd194: data = 1'd1;
		12'd195: data = 1'd1;
		12'd196: data = 1'd1;
		12'd197: data = 1'd1;
		12'd198: data = 1'd1;
		12'd199: data = 1'd0;
		12'd200: data = 1'd1;
		12'd201: data = 1'd1;
		12'd202: data = 1'd1;
		12'd203: data = 1'd1;
		12'd204: data = 1'd1;
		12'd205: data = 1'd1;
		12'd206: data = 1'd1;
		12'd207: data = 1'd1;
		12'd208: data = 1'd0;
		12'd209: data = 1'd0;
		12'd210: data = 1'd0;
		12'd211: data = 1'd0;
		12'd212: data = 1'd0;
		12'd213: data = 1'd0;
		12'd214: data = 1'd1;
		12'd215: data = 1'd0;
		12'd216: data = 1'd1;
		12'd217: data = 1'd1;
		12'd218: data = 1'd1;
		12'd219: data = 1'd1;
		12'd220: data = 1'd1;
		12'd221: data = 1'd1;
		12'd222: data = 1'd1;
		12'd223: data = 1'd1;
		12'd224: data = 1'd1;
		12'd225: data = 1'd1;
		12'd226: data = 1'd1;
		12'd227: data = 1'd1;
		12'd228: data = 1'd1;
		12'd229: data = 1'd0;
		12'd230: data = 1'd1;
		12'd231: data = 1'd1;
		12'd232: data = 1'd0;
		12'd233: data = 1'd1;
		12'd234: data = 1'd1;
		12'd235: data = 1'd1;
		12'd236: data = 1'd1;
		12'd237: data = 1'd1;
		12'd238: data = 1'd1;
		12'd239: data = 1'd1;
		12'd240: data = 1'd1;
		12'd241: data = 1'd0;
		12'd242: data = 1'd0;
		12'd243: data = 1'd0;
		12'd244: data = 1'd0;
		12'd245: data = 1'd1;
		12'd246: data = 1'd0;
		12'd247: data = 1'd1;
		12'd248: data = 1'd0;
		12'd249: data = 1'd1;
		12'd250: data = 1'd1;
		12'd251: data = 1'd1;
		12'd252: data = 1'd1;
		12'd253: data = 1'd1;
		12'd254: data = 1'd1;
		12'd255: data = 1'd1;
		12'd256: data = 1'd1;
		12'd257: data = 1'd0;
		12'd258: data = 1'd0;
		12'd259: data = 1'd0;
		12'd260: data = 1'd0;
		12'd261: data = 1'd0;
		12'd262: data = 1'd1;
		12'd263: data = 1'd0;
		12'd264: data = 1'd1;
		12'd265: data = 1'd1;
		12'd266: data = 1'd1;
		12'd267: data = 1'd1;
		12'd268: data = 1'd1;
		12'd269: data = 1'd1;
		12'd270: data = 1'd1;
		12'd271: data = 1'd1;
		12'd272: data = 1'd1;
		12'd273: data = 1'd1;
		12'd274: data = 1'd1;
		12'd275: data = 1'd1;
		12'd276: data = 1'd1;
		12'd277: data = 1'd1;
		12'd278: data = 1'd1;
		12'd279: data = 1'd1;
		12'd280: data = 1'd0;
		12'd281: data = 1'd1;
		12'd282: data = 1'd1;
		12'd283: data = 1'd1;
		12'd284: data = 1'd1;
		12'd285: data = 1'd1;
		12'd286: data = 1'd1;
		12'd287: data = 1'd1;
		12'd288: data = 1'd1;
		12'd289: data = 1'd1;
		12'd290: data = 1'd1;
		12'd291: data = 1'd1;
		12'd292: data = 1'd1;
		12'd293: data = 1'd1;
		12'd294: data = 1'd1;
		12'd295: data = 1'd1;
		12'd296: data = 1'd1;
		12'd297: data = 1'd0;
		12'd298: data = 1'd0;
		12'd299: data = 1'd1;
		12'd300: data = 1'd1;
		12'd301: data = 1'd1;
		12'd302: data = 1'd1;
		12'd303: data = 1'd1;
		12'd304: data = 1'd1;
		12'd305: data = 1'd1;
		12'd306: data = 1'd1;
		12'd307: data = 1'd1;
		12'd308: data = 1'd1;
		12'd309: data = 1'd1;
		12'd310: data = 1'd1;
		12'd311: data = 1'd1;
		12'd312: data = 1'd1;
		12'd313: data = 1'd1;
		12'd314: data = 1'd0;
		12'd315: data = 1'd0;
		12'd316: data = 1'd1;
		12'd317: data = 1'd1;
		12'd318: data = 1'd1;
		12'd319: data = 1'd1;
		12'd320: data = 1'd1;
		12'd321: data = 1'd1;
		12'd322: data = 1'd1;
		12'd323: data = 1'd1;
		12'd324: data = 1'd1;
		12'd325: data = 1'd1;
		12'd326: data = 1'd1;
		12'd327: data = 1'd1;
		12'd328: data = 1'd1;
		12'd329: data = 1'd1;
		12'd330: data = 1'd0;
		12'd331: data = 1'd0;
		12'd332: data = 1'd0;
		12'd333: data = 1'd1;
		12'd334: data = 1'd1;
		12'd335: data = 1'd1;
		12'd336: data = 1'd1;
		12'd337: data = 1'd1;
		12'd338: data = 1'd1;
		12'd339: data = 1'd1;
		12'd340: data = 1'd1;
		12'd341: data = 1'd1;
		12'd342: data = 1'd1;
		12'd343: data = 1'd1;
		12'd344: data = 1'd1;
		12'd345: data = 1'd0;
		12'd346: data = 1'd0;
		12'd347: data = 1'd0;
		12'd348: data = 1'd0;
		12'd349: data = 1'd1;
		12'd350: data = 1'd1;
		12'd351: data = 1'd1;
		12'd352: data = 1'd0;
		12'd353: data = 1'd1;
		12'd354: data = 1'd1;
		12'd355: data = 1'd1;
		12'd356: data = 1'd1;
		12'd357: data = 1'd1;
		12'd358: data = 1'd1;
		12'd359: data = 1'd0;
		12'd360: data = 1'd0;
		12'd361: data = 1'd0;
		12'd362: data = 1'd0;
		12'd363: data = 1'd1;
		12'd364: data = 1'd1;
		12'd365: data = 1'd1;
		12'd366: data = 1'd1;
		12'd367: data = 1'd1;
		12'd368: data = 1'd0;
		12'd369: data = 1'd0;
		12'd370: data = 1'd1;
		12'd371: data = 1'd1;
		12'd372: data = 1'd1;
		12'd373: data = 1'd1;
		12'd374: data = 1'd1;
		12'd375: data = 1'd1;
		12'd376: data = 1'd0;
		12'd377: data = 1'd1;
		12'd378: data = 1'd1;
		12'd379: data = 1'd1;
		12'd380: data = 1'd1;
		12'd381: data = 1'd1;
		12'd382: data = 1'd1;
		12'd383: data = 1'd1;
		12'd384: data = 1'd0;
		12'd385: data = 1'd0;
		12'd386: data = 1'd0;
		12'd387: data = 1'd1;
		12'd388: data = 1'd1;
		12'd389: data = 1'd1;
		12'd390: data = 1'd1;
		12'd391: data = 1'd1;
		12'd392: data = 1'd0;
		12'd393: data = 1'd1;
		12'd394: data = 1'd1;
		12'd395: data = 1'd1;
		12'd396: data = 1'd1;
		12'd397: data = 1'd1;
		12'd398: data = 1'd1;
		12'd399: data = 1'd1;
		12'd400: data = 1'd0;
		12'd401: data = 1'd0;
		12'd402: data = 1'd0;
		12'd403: data = 1'd0;
		12'd404: data = 1'd1;
		12'd405: data = 1'd1;
		12'd406: data = 1'd1;
		12'd407: data = 1'd1;
		12'd408: data = 1'd0;
		12'd409: data = 1'd1;
		12'd410: data = 1'd1;
		12'd411: data = 1'd1;
		12'd412: data = 1'd1;
		12'd413: data = 1'd1;
		12'd414: data = 1'd1;
		12'd415: data = 1'd1;
		12'd416: data = 1'd0;
		12'd417: data = 1'd0;
		12'd418: data = 1'd0;
		12'd419: data = 1'd0;
		12'd420: data = 1'd1;
		12'd421: data = 1'd1;
		12'd422: data = 1'd1;
		12'd423: data = 1'd1;
		12'd424: data = 1'd0;
		12'd425: data = 1'd1;
		12'd426: data = 1'd1;
		12'd427: data = 1'd1;
		12'd428: data = 1'd1;
		12'd429: data = 1'd1;
		12'd430: data = 1'd1;
		12'd431: data = 1'd1;
		12'd432: data = 1'd0;
		12'd433: data = 1'd0;
		12'd434: data = 1'd0;
		12'd435: data = 1'd0;
		12'd436: data = 1'd0;
		12'd437: data = 1'd0;
		12'd438: data = 1'd0;
		12'd439: data = 1'd1;
		12'd440: data = 1'd0;
		12'd441: data = 1'd1;
		12'd442: data = 1'd1;
		12'd443: data = 1'd1;
		12'd444: data = 1'd1;
		12'd445: data = 1'd1;
		12'd446: data = 1'd1;
		12'd447: data = 1'd1;
		12'd448: data = 1'd1;
		12'd449: data = 1'd1;
		12'd450: data = 1'd1;
		12'd451: data = 1'd1;
		12'd452: data = 1'd1;
		12'd453: data = 1'd1;
		12'd454: data = 1'd0;
		12'd455: data = 1'd1;
		12'd456: data = 1'd1;
		12'd457: data = 1'd0;
		12'd458: data = 1'd1;
		12'd459: data = 1'd1;
		12'd460: data = 1'd1;
		12'd461: data = 1'd1;
		12'd462: data = 1'd1;
		12'd463: data = 1'd1;
		12'd464: data = 1'd0;
		12'd465: data = 1'd0;
		12'd466: data = 1'd0;
		12'd467: data = 1'd0;
		12'd468: data = 1'd0;
		12'd469: data = 1'd0;
		12'd470: data = 1'd1;
		12'd471: data = 1'd0;
		12'd472: data = 1'd1;
		12'd473: data = 1'd0;
		12'd474: data = 1'd1;
		12'd475: data = 1'd1;
		12'd476: data = 1'd1;
		12'd477: data = 1'd1;
		12'd478: data = 1'd1;
		12'd479: data = 1'd1;
		12'd480: data = 1'd1;
		12'd481: data = 1'd0;
		12'd482: data = 1'd1;
		12'd483: data = 1'd1;
		12'd484: data = 1'd1;
		12'd485: data = 1'd0;
		12'd486: data = 1'd1;
		12'd487: data = 1'd0;
		12'd488: data = 1'd1;
		12'd489: data = 1'd0;
		12'd490: data = 1'd0;
		12'd491: data = 1'd1;
		12'd492: data = 1'd1;
		12'd493: data = 1'd1;
		12'd494: data = 1'd1;
		12'd495: data = 1'd1;
		12'd496: data = 1'd1;
		12'd497: data = 1'd0;
		12'd498: data = 1'd1;
		12'd499: data = 1'd0;
		12'd500: data = 1'd1;
		12'd501: data = 1'd0;
		12'd502: data = 1'd1;
		12'd503: data = 1'd1;
		12'd504: data = 1'd0;
		12'd505: data = 1'd1;
		12'd506: data = 1'd0;
		12'd507: data = 1'd1;
		12'd508: data = 1'd1;
		12'd509: data = 1'd1;
		12'd510: data = 1'd1;
		12'd511: data = 1'd1;
		12'd512: data = 1'd1;
		12'd513: data = 1'd1;
		12'd514: data = 1'd0;
		12'd515: data = 1'd0;
		12'd516: data = 1'd0;
		12'd517: data = 1'd0;
		12'd518: data = 1'd0;
		12'd519: data = 1'd0;
		12'd520: data = 1'd1;
		12'd521: data = 1'd0;
		12'd522: data = 1'd0;
		12'd523: data = 1'd1;
		12'd524: data = 1'd1;
		12'd525: data = 1'd1;
		12'd526: data = 1'd1;
		12'd527: data = 1'd1;
		12'd528: data = 1'd1;
		12'd529: data = 1'd0;
		12'd530: data = 1'd0;
		12'd531: data = 1'd0;
		12'd532: data = 1'd0;
		12'd533: data = 1'd0;
		12'd534: data = 1'd1;
		12'd535: data = 1'd0;
		12'd536: data = 1'd1;
		12'd537: data = 1'd1;
		12'd538: data = 1'd0;
		12'd539: data = 1'd0;
		12'd540: data = 1'd1;
		12'd541: data = 1'd1;
		12'd542: data = 1'd1;
		12'd543: data = 1'd1;
		12'd544: data = 1'd1;
		12'd545: data = 1'd0;
		12'd546: data = 1'd0;
		12'd547: data = 1'd0;
		12'd548: data = 1'd0;
		12'd549: data = 1'd0;
		12'd550: data = 1'd0;
		12'd551: data = 1'd1;
		12'd552: data = 1'd0;
		12'd553: data = 1'd1;
		12'd554: data = 1'd1;
		12'd555: data = 1'd0;
		12'd556: data = 1'd0;
		12'd557: data = 1'd1;
		12'd558: data = 1'd1;
		12'd559: data = 1'd1;
		12'd560: data = 1'd1;
		12'd561: data = 1'd0;
		12'd562: data = 1'd0;
		12'd563: data = 1'd0;
		12'd564: data = 1'd0;
		12'd565: data = 1'd0;
		12'd566: data = 1'd0;
		12'd567: data = 1'd0;
		12'd568: data = 1'd1;
		12'd569: data = 1'd0;
		12'd570: data = 1'd1;
		12'd571: data = 1'd1;
		12'd572: data = 1'd0;
		12'd573: data = 1'd0;
		12'd574: data = 1'd0;
		12'd575: data = 1'd1;
		12'd576: data = 1'd1;
		12'd577: data = 1'd0;
		12'd578: data = 1'd0;
		12'd579: data = 1'd0;
		12'd580: data = 1'd0;
		12'd581: data = 1'd0;
		12'd582: data = 1'd0;
		12'd583: data = 1'd0;
		12'd584: data = 1'd1;
		12'd585: data = 1'd0;
		12'd586: data = 1'd0;
		12'd587: data = 1'd1;
		12'd588: data = 1'd1;
		12'd589: data = 1'd1;
		12'd590: data = 1'd0;
		12'd591: data = 1'd0;
		12'd592: data = 1'd1;
		12'd593: data = 1'd1;
		12'd594: data = 1'd1;
		12'd595: data = 1'd1;
		12'd596: data = 1'd1;
		12'd597: data = 1'd1;
		12'd598: data = 1'd1;
		12'd599: data = 1'd1;
		12'd600: data = 1'd1;
		12'd601: data = 1'd0;
		12'd602: data = 1'd0;
		12'd603: data = 1'd0;
		12'd604: data = 1'd1;
		12'd605: data = 1'd1;
		12'd606: data = 1'd1;
		12'd607: data = 1'd0;
		12'd608: data = 1'd1;
		12'd609: data = 1'd1;
		12'd610: data = 1'd1;
		12'd611: data = 1'd1;
		12'd612: data = 1'd1;
		12'd613: data = 1'd1;
		12'd614: data = 1'd1;
		12'd615: data = 1'd1;
		12'd616: data = 1'd0;
		12'd617: data = 1'd0;
		12'd618: data = 1'd0;
		12'd619: data = 1'd1;
		12'd620: data = 1'd1;
		12'd621: data = 1'd1;
		12'd622: data = 1'd1;
		12'd623: data = 1'd0;
		12'd624: data = 1'd0;
		12'd625: data = 1'd0;
		12'd626: data = 1'd1;
		12'd627: data = 1'd1;
		12'd628: data = 1'd1;
		12'd629: data = 1'd1;
		12'd630: data = 1'd1;
		12'd631: data = 1'd1;
		12'd632: data = 1'd0;
		12'd633: data = 1'd1;
		12'd634: data = 1'd1;
		12'd635: data = 1'd1;
		12'd636: data = 1'd1;
		12'd637: data = 1'd1;
		12'd638: data = 1'd0;
		12'd639: data = 1'd0;
		12'd640: data = 1'd0;
		12'd641: data = 1'd0;
		12'd642: data = 1'd0;
		12'd643: data = 1'd1;
		12'd644: data = 1'd1;
		12'd645: data = 1'd1;
		12'd646: data = 1'd1;
		12'd647: data = 1'd1;
		12'd648: data = 1'd0;
		12'd649: data = 1'd1;
		12'd650: data = 1'd0;
		12'd651: data = 1'd1;
		12'd652: data = 1'd0;
		12'd653: data = 1'd0;
		12'd654: data = 1'd0;
		12'd655: data = 1'd0;
		12'd656: data = 1'd0;
		12'd657: data = 1'd0;
		12'd658: data = 1'd0;
		12'd659: data = 1'd1;
		12'd660: data = 1'd1;
		12'd661: data = 1'd1;
		12'd662: data = 1'd1;
		12'd663: data = 1'd1;
		12'd664: data = 1'd0;
		12'd665: data = 1'd1;
		12'd666: data = 1'd0;
		12'd667: data = 1'd0;
		12'd668: data = 1'd0;
		12'd669: data = 1'd0;
		12'd670: data = 1'd0;
		12'd671: data = 1'd0;
		12'd672: data = 1'd0;
		12'd673: data = 1'd0;
		12'd674: data = 1'd0;
		12'd675: data = 1'd0;
		12'd676: data = 1'd1;
		12'd677: data = 1'd1;
		12'd678: data = 1'd1;
		12'd679: data = 1'd1;
		12'd680: data = 1'd0;
		12'd681: data = 1'd1;
		12'd682: data = 1'd0;
		12'd683: data = 1'd1;
		12'd684: data = 1'd1;
		12'd685: data = 1'd0;
		12'd686: data = 1'd0;
		12'd687: data = 1'd0;
		12'd688: data = 1'd0;
		12'd689: data = 1'd0;
		12'd690: data = 1'd0;
		12'd691: data = 1'd0;
		12'd692: data = 1'd0;
		12'd693: data = 1'd0;
		12'd694: data = 1'd0;
		12'd695: data = 1'd1;
		12'd696: data = 1'd0;
		12'd697: data = 1'd1;
		12'd698: data = 1'd0;
		12'd699: data = 1'd1;
		12'd700: data = 1'd1;
		12'd701: data = 1'd1;
		12'd702: data = 1'd1;
		12'd703: data = 1'd1;
		12'd704: data = 1'd0;
		12'd705: data = 1'd1;
		12'd706: data = 1'd1;
		12'd707: data = 1'd1;
		12'd708: data = 1'd1;
		12'd709: data = 1'd1;
		12'd710: data = 1'd0;
		12'd711: data = 1'd1;
		12'd712: data = 1'd0;
		12'd713: data = 1'd1;
		12'd714: data = 1'd0;
		12'd715: data = 1'd0;
		12'd716: data = 1'd1;
		12'd717: data = 1'd1;
		12'd718: data = 1'd1;
		12'd719: data = 1'd1;
		12'd720: data = 1'd0;
		12'd721: data = 1'd1;
		12'd722: data = 1'd1;
		12'd723: data = 1'd0;
		12'd724: data = 1'd1;
		12'd725: data = 1'd1;
		12'd726: data = 1'd0;
		12'd727: data = 1'd1;
		12'd728: data = 1'd1;
		12'd729: data = 1'd0;
		12'd730: data = 1'd1;
		12'd731: data = 1'd0;
		12'd732: data = 1'd1;
		12'd733: data = 1'd1;
		12'd734: data = 1'd1;
		12'd735: data = 1'd1;
		12'd736: data = 1'd0;
		12'd737: data = 1'd0;
		12'd738: data = 1'd1;
		12'd739: data = 1'd0;
		12'd740: data = 1'd1;
		12'd741: data = 1'd0;
		12'd742: data = 1'd1;
		12'd743: data = 1'd0;
		12'd744: data = 1'd1;
		12'd745: data = 1'd0;
		12'd746: data = 1'd1;
		12'd747: data = 1'd0;
		12'd748: data = 1'd1;
		12'd749: data = 1'd1;
		12'd750: data = 1'd1;
		12'd751: data = 1'd1;
		12'd752: data = 1'd1;
		12'd753: data = 1'd0;
		12'd754: data = 1'd1;
		12'd755: data = 1'd0;
		12'd756: data = 1'd1;
		12'd757: data = 1'd1;
		12'd758: data = 1'd0;
		12'd759: data = 1'd0;
		12'd760: data = 1'd1;
		12'd761: data = 1'd0;
		12'd762: data = 1'd0;
		12'd763: data = 1'd1;
		12'd764: data = 1'd0;
		12'd765: data = 1'd1;
		12'd766: data = 1'd1;
		12'd767: data = 1'd1;
		12'd768: data = 1'd1;
		12'd769: data = 1'd0;
		12'd770: data = 1'd0;
		12'd771: data = 1'd0;
		12'd772: data = 1'd0;
		12'd773: data = 1'd1;
		12'd774: data = 1'd0;
		12'd775: data = 1'd1;
		12'd776: data = 1'd0;
		12'd777: data = 1'd1;
		12'd778: data = 1'd1;
		12'd779: data = 1'd0;
		12'd780: data = 1'd0;
		12'd781: data = 1'd0;
		12'd782: data = 1'd0;
		12'd783: data = 1'd1;
		12'd784: data = 1'd1;
		12'd785: data = 1'd1;
		12'd786: data = 1'd1;
		12'd787: data = 1'd1;
		12'd788: data = 1'd1;
		12'd789: data = 1'd1;
		12'd790: data = 1'd0;
		12'd791: data = 1'd1;
		12'd792: data = 1'd0;
		12'd793: data = 1'd0;
		12'd794: data = 1'd1;
		12'd795: data = 1'd1;
		12'd796: data = 1'd1;
		12'd797: data = 1'd0;
		12'd798: data = 1'd0;
		12'd799: data = 1'd0;
		12'd800: data = 1'd1;
		12'd801: data = 1'd1;
		12'd802: data = 1'd1;
		12'd803: data = 1'd1;
		12'd804: data = 1'd1;
		12'd805: data = 1'd0;
		12'd806: data = 1'd1;
		12'd807: data = 1'd0;
		12'd808: data = 1'd1;
		12'd809: data = 1'd0;
		12'd810: data = 1'd0;
		12'd811: data = 1'd0;
		12'd812: data = 1'd1;
		12'd813: data = 1'd1;
		12'd814: data = 1'd0;
		12'd815: data = 1'd0;
		12'd816: data = 1'd1;
		12'd817: data = 1'd1;
		12'd818: data = 1'd1;
		12'd819: data = 1'd1;
		12'd820: data = 1'd1;
		12'd821: data = 1'd1;
		12'd822: data = 1'd0;
		12'd823: data = 1'd1;
		12'd824: data = 1'd0;
		12'd825: data = 1'd1;
		12'd826: data = 1'd0;
		12'd827: data = 1'd0;
		12'd828: data = 1'd0;
		12'd829: data = 1'd1;
		12'd830: data = 1'd1;
		12'd831: data = 1'd0;
		12'd832: data = 1'd1;
		12'd833: data = 1'd0;
		12'd834: data = 1'd0;
		12'd835: data = 1'd0;
		12'd836: data = 1'd0;
		12'd837: data = 1'd0;
		12'd838: data = 1'd0;
		12'd839: data = 1'd1;
		12'd840: data = 1'd1;
		12'd841: data = 1'd0;
		12'd842: data = 1'd1;
		12'd843: data = 1'd1;
		12'd844: data = 1'd0;
		12'd845: data = 1'd0;
		12'd846: data = 1'd1;
		12'd847: data = 1'd1;
		12'd848: data = 1'd1;
		12'd849: data = 1'd0;
		12'd850: data = 1'd0;
		12'd851: data = 1'd0;
		12'd852: data = 1'd0;
		12'd853: data = 1'd0;
		12'd854: data = 1'd0;
		12'd855: data = 1'd0;
		12'd856: data = 1'd1;
		12'd857: data = 1'd0;
		12'd858: data = 1'd0;
		12'd859: data = 1'd1;
		12'd860: data = 1'd1;
		12'd861: data = 1'd0;
		12'd862: data = 1'd0;
		12'd863: data = 1'd1;
		12'd864: data = 1'd1;
		12'd865: data = 1'd0;
		12'd866: data = 1'd0;
		12'd867: data = 1'd0;
		12'd868: data = 1'd0;
		12'd869: data = 1'd0;
		12'd870: data = 1'd0;
		12'd871: data = 1'd1;
		12'd872: data = 1'd0;
		12'd873: data = 1'd0;
		12'd874: data = 1'd1;
		12'd875: data = 1'd1;
		12'd876: data = 1'd1;
		12'd877: data = 1'd1;
		12'd878: data = 1'd0;
		12'd879: data = 1'd0;
		12'd880: data = 1'd1;
		12'd881: data = 1'd0;
		12'd882: data = 1'd0;
		12'd883: data = 1'd0;
		12'd884: data = 1'd0;
		12'd885: data = 1'd0;
		12'd886: data = 1'd0;
		12'd887: data = 1'd1;
		12'd888: data = 1'd0;
		12'd889: data = 1'd1;
		12'd890: data = 1'd1;
		12'd891: data = 1'd1;
		12'd892: data = 1'd1;
		12'd893: data = 1'd0;
		12'd894: data = 1'd0;
		12'd895: data = 1'd0;
		12'd896: data = 1'd1;
		12'd897: data = 1'd0;
		12'd898: data = 1'd0;
		12'd899: data = 1'd0;
		12'd900: data = 1'd0;
		12'd901: data = 1'd0;
		12'd902: data = 1'd0;
		12'd903: data = 1'd1;
		12'd904: data = 1'd0;
		12'd905: data = 1'd1;
		12'd906: data = 1'd1;
		12'd907: data = 1'd1;
		12'd908: data = 1'd0;
		12'd909: data = 1'd0;
		12'd910: data = 1'd0;
		12'd911: data = 1'd0;
		12'd912: data = 1'd0;
		12'd913: data = 1'd0;
		12'd914: data = 1'd0;
		12'd915: data = 1'd1;
		12'd916: data = 1'd1;
		12'd917: data = 1'd1;
		12'd918: data = 1'd1;
		12'd919: data = 1'd1;
		12'd920: data = 1'd0;
		12'd921: data = 1'd1;
		12'd922: data = 1'd0;
		12'd923: data = 1'd0;
		12'd924: data = 1'd0;
		12'd925: data = 1'd0;
		12'd926: data = 1'd0;
		12'd927: data = 1'd1;
		12'd928: data = 1'd1;
		12'd929: data = 1'd0;
		12'd930: data = 1'd0;
		12'd931: data = 1'd0;
		12'd932: data = 1'd1;
		12'd933: data = 1'd1;
		12'd934: data = 1'd1;
		12'd935: data = 1'd0;
		12'd936: data = 1'd1;
		12'd937: data = 1'd0;
		12'd938: data = 1'd1;
		12'd939: data = 1'd1;
		12'd940: data = 1'd0;
		12'd941: data = 1'd0;
		12'd942: data = 1'd1;
		12'd943: data = 1'd1;
		12'd944: data = 1'd0;
		12'd945: data = 1'd1;
		12'd946: data = 1'd0;
		12'd947: data = 1'd0;
		12'd948: data = 1'd0;
		12'd949: data = 1'd1;
		12'd950: data = 1'd1;
		12'd951: data = 1'd0;
		12'd952: data = 1'd1;
		12'd953: data = 1'd1;
		12'd954: data = 1'd0;
		12'd955: data = 1'd1;
		12'd956: data = 1'd0;
		12'd957: data = 1'd1;
		12'd958: data = 1'd1;
		12'd959: data = 1'd1;
		12'd960: data = 1'd0;
		12'd961: data = 1'd1;
		12'd962: data = 1'd0;
		12'd963: data = 1'd1;
		12'd964: data = 1'd1;
		12'd965: data = 1'd0;
		12'd966: data = 1'd0;
		12'd967: data = 1'd1;
		12'd968: data = 1'd0;
		12'd969: data = 1'd1;
		12'd970: data = 1'd0;
		12'd971: data = 1'd1;
		12'd972: data = 1'd0;
		12'd973: data = 1'd0;
		12'd974: data = 1'd0;
		12'd975: data = 1'd0;
		12'd976: data = 1'd0;
		12'd977: data = 1'd1;
		12'd978: data = 1'd0;
		12'd979: data = 1'd0;
		12'd980: data = 1'd1;
		12'd981: data = 1'd0;
		12'd982: data = 1'd0;
		12'd983: data = 1'd1;
		12'd984: data = 1'd0;
		12'd985: data = 1'd1;
		12'd986: data = 1'd0;
		12'd987: data = 1'd0;
		12'd988: data = 1'd1;
		12'd989: data = 1'd0;
		12'd990: data = 1'd1;
		12'd991: data = 1'd1;
		12'd992: data = 1'd0;
		12'd993: data = 1'd0;
		12'd994: data = 1'd1;
		12'd995: data = 1'd0;
		12'd996: data = 1'd1;
		12'd997: data = 1'd1;
		12'd998: data = 1'd0;
		12'd999: data = 1'd0;
		12'd1000: data = 1'd1;
		12'd1001: data = 1'd0;
		12'd1002: data = 1'd1;
		12'd1003: data = 1'd0;
		12'd1004: data = 1'd1;
		12'd1005: data = 1'd0;
		12'd1006: data = 1'd1;
		12'd1007: data = 1'd1;
		12'd1008: data = 1'd0;
		12'd1009: data = 1'd0;
		12'd1010: data = 1'd0;
		12'd1011: data = 1'd0;
		12'd1012: data = 1'd1;
		12'd1013: data = 1'd1;
		12'd1014: data = 1'd0;
		12'd1015: data = 1'd0;
		12'd1016: data = 1'd0;
		12'd1017: data = 1'd1;
		12'd1018: data = 1'd1;
		12'd1019: data = 1'd0;
		12'd1020: data = 1'd1;
		12'd1021: data = 1'd1;
		12'd1022: data = 1'd0;
		12'd1023: data = 1'd1;
		12'd1024: data = 1'd1;
		12'd1025: data = 1'd0;
		12'd1026: data = 1'd1;
		12'd1027: data = 1'd0;
		12'd1028: data = 1'd1;
		12'd1029: data = 1'd1;
		12'd1030: data = 1'd0;
		12'd1031: data = 1'd1;
		12'd1032: data = 1'd0;
		12'd1033: data = 1'd1;
		12'd1034: data = 1'd1;
		12'd1035: data = 1'd0;
		12'd1036: data = 1'd0;
		12'd1037: data = 1'd1;
		12'd1038: data = 1'd1;
		12'd1039: data = 1'd1;
		12'd1040: data = 1'd1;
		12'd1041: data = 1'd0;
		12'd1042: data = 1'd1;
		12'd1043: data = 1'd0;
		12'd1044: data = 1'd0;
		12'd1045: data = 1'd1;
		12'd1046: data = 1'd0;
		12'd1047: data = 1'd1;
		12'd1048: data = 1'd0;
		12'd1049: data = 1'd1;
		12'd1050: data = 1'd1;
		12'd1051: data = 1'd0;
		12'd1052: data = 1'd0;
		12'd1053: data = 1'd0;
		12'd1054: data = 1'd1;
		12'd1055: data = 1'd1;
		12'd1056: data = 1'd1;
		12'd1057: data = 1'd1;
		12'd1058: data = 1'd0;
		12'd1059: data = 1'd0;
		12'd1060: data = 1'd0;
		12'd1061: data = 1'd1;
		12'd1062: data = 1'd0;
		12'd1063: data = 1'd1;
		12'd1064: data = 1'd0;
		12'd1065: data = 1'd0;
		12'd1066: data = 1'd1;
		12'd1067: data = 1'd1;
		12'd1068: data = 1'd0;
		12'd1069: data = 1'd0;
		12'd1070: data = 1'd0;
		12'd1071: data = 1'd1;
		12'd1072: data = 1'd1;
		12'd1073: data = 1'd1;
		12'd1074: data = 1'd1;
		12'd1075: data = 1'd1;
		12'd1076: data = 1'd1;
		12'd1077: data = 1'd0;
		12'd1078: data = 1'd1;
		12'd1079: data = 1'd0;
		12'd1080: data = 1'd1;
		12'd1081: data = 1'd0;
		12'd1082: data = 1'd0;
		12'd1083: data = 1'd1;
		12'd1084: data = 1'd1;
		12'd1085: data = 1'd1;
		12'd1086: data = 1'd0;
		12'd1087: data = 1'd0;
		12'd1088: data = 1'd1;
		12'd1089: data = 1'd1;
		12'd1090: data = 1'd1;
		12'd1091: data = 1'd1;
		12'd1092: data = 1'd1;
		12'd1093: data = 1'd1;
		12'd1094: data = 1'd0;
		12'd1095: data = 1'd1;
		12'd1096: data = 1'd0;
		12'd1097: data = 1'd1;
		12'd1098: data = 1'd0;
		12'd1099: data = 1'd0;
		12'd1100: data = 1'd1;
		12'd1101: data = 1'd1;
		12'd1102: data = 1'd1;
		12'd1103: data = 1'd0;
		12'd1104: data = 1'd1;
		12'd1105: data = 1'd1;
		12'd1106: data = 1'd1;
		12'd1107: data = 1'd1;
		12'd1108: data = 1'd1;
		12'd1109: data = 1'd1;
		12'd1110: data = 1'd0;
		12'd1111: data = 1'd1;
		12'd1112: data = 1'd0;
		12'd1113: data = 1'd1;
		12'd1114: data = 1'd1;
		12'd1115: data = 1'd0;
		12'd1116: data = 1'd0;
		12'd1117: data = 1'd0;
		12'd1118: data = 1'd1;
		12'd1119: data = 1'd1;
		12'd1120: data = 1'd1;
		12'd1121: data = 1'd1;
		12'd1122: data = 1'd1;
		12'd1123: data = 1'd1;
		12'd1124: data = 1'd1;
		12'd1125: data = 1'd1;
		12'd1126: data = 1'd0;
		12'd1127: data = 1'd1;
		12'd1128: data = 1'd0;
		12'd1129: data = 1'd0;
		12'd1130: data = 1'd1;
		12'd1131: data = 1'd1;
		12'd1132: data = 1'd0;
		12'd1133: data = 1'd0;
		12'd1134: data = 1'd0;
		12'd1135: data = 1'd1;
		12'd1136: data = 1'd1;
		12'd1137: data = 1'd1;
		12'd1138: data = 1'd1;
		12'd1139: data = 1'd1;
		12'd1140: data = 1'd1;
		12'd1141: data = 1'd1;
		12'd1142: data = 1'd0;
		12'd1143: data = 1'd1;
		12'd1144: data = 1'd0;
		12'd1145: data = 1'd0;
		12'd1146: data = 1'd1;
		12'd1147: data = 1'd1;
		12'd1148: data = 1'd1;
		12'd1149: data = 1'd0;
		12'd1150: data = 1'd0;
		12'd1151: data = 1'd0;
		12'd1152: data = 1'd1;
		12'd1153: data = 1'd0;
		12'd1154: data = 1'd0;
		12'd1155: data = 1'd0;
		12'd1156: data = 1'd0;
		12'd1157: data = 1'd0;
		12'd1158: data = 1'd0;
		12'd1159: data = 1'd1;
		12'd1160: data = 1'd0;
		12'd1161: data = 1'd1;
		12'd1162: data = 1'd1;
		12'd1163: data = 1'd1;
		12'd1164: data = 1'd0;
		12'd1165: data = 1'd0;
		12'd1166: data = 1'd0;
		12'd1167: data = 1'd0;
		12'd1168: data = 1'd1;
		12'd1169: data = 1'd1;
		12'd1170: data = 1'd0;
		12'd1171: data = 1'd0;
		12'd1172: data = 1'd0;
		12'd1173: data = 1'd0;
		12'd1174: data = 1'd1;
		12'd1175: data = 1'd1;
		12'd1176: data = 1'd0;
		12'd1177: data = 1'd1;
		12'd1178: data = 1'd1;
		12'd1179: data = 1'd0;
		12'd1180: data = 1'd0;
		12'd1181: data = 1'd0;
		12'd1182: data = 1'd0;
		12'd1183: data = 1'd0;
		12'd1184: data = 1'd0;
		12'd1185: data = 1'd0;
		12'd1186: data = 1'd1;
		12'd1187: data = 1'd0;
		12'd1188: data = 1'd0;
		12'd1189: data = 1'd0;
		12'd1190: data = 1'd1;
		12'd1191: data = 1'd1;
		12'd1192: data = 1'd0;
		12'd1193: data = 1'd1;
		12'd1194: data = 1'd1;
		12'd1195: data = 1'd0;
		12'd1196: data = 1'd0;
		12'd1197: data = 1'd0;
		12'd1198: data = 1'd0;
		12'd1199: data = 1'd1;
		12'd1200: data = 1'd0;
		12'd1201: data = 1'd1;
		12'd1202: data = 1'd0;
		12'd1203: data = 1'd1;
		12'd1204: data = 1'd1;
		12'd1205: data = 1'd0;
		12'd1206: data = 1'd1;
		12'd1207: data = 1'd1;
		12'd1208: data = 1'd0;
		12'd1209: data = 1'd1;
		12'd1210: data = 1'd1;
		12'd1211: data = 1'd0;
		12'd1212: data = 1'd1;
		12'd1213: data = 1'd0;
		12'd1214: data = 1'd1;
		12'd1215: data = 1'd1;
		12'd1216: data = 1'd0;
		12'd1217: data = 1'd1;
		12'd1218: data = 1'd0;
		12'd1219: data = 1'd1;
		12'd1220: data = 1'd0;
		12'd1221: data = 1'd0;
		12'd1222: data = 1'd0;
		12'd1223: data = 1'd1;
		12'd1224: data = 1'd0;
		12'd1225: data = 1'd1;
		12'd1226: data = 1'd1;
		12'd1227: data = 1'd0;
		12'd1228: data = 1'd1;
		12'd1229: data = 1'd1;
		12'd1230: data = 1'd1;
		12'd1231: data = 1'd1;
		12'd1232: data = 1'd0;
		12'd1233: data = 1'd0;
		12'd1234: data = 1'd0;
		12'd1235: data = 1'd0;
		12'd1236: data = 1'd1;
		12'd1237: data = 1'd0;
		12'd1238: data = 1'd0;
		12'd1239: data = 1'd0;
		12'd1240: data = 1'd1;
		12'd1241: data = 1'd1;
		12'd1242: data = 1'd1;
		12'd1243: data = 1'd0;
		12'd1244: data = 1'd1;
		12'd1245: data = 1'd1;
		12'd1246: data = 1'd0;
		12'd1247: data = 1'd0;
		12'd1248: data = 1'd0;
		12'd1249: data = 1'd0;
		12'd1250: data = 1'd0;
		12'd1251: data = 1'd0;
		12'd1252: data = 1'd0;
		12'd1253: data = 1'd1;
		12'd1254: data = 1'd0;
		12'd1255: data = 1'd0;
		12'd1256: data = 1'd0;
		12'd1257: data = 1'd1;
		12'd1258: data = 1'd1;
		12'd1259: data = 1'd0;
		12'd1260: data = 1'd1;
		12'd1261: data = 1'd1;
		12'd1262: data = 1'd0;
		12'd1263: data = 1'd1;
		12'd1264: data = 1'd0;
		12'd1265: data = 1'd0;
		12'd1266: data = 1'd0;
		12'd1267: data = 1'd0;
		12'd1268: data = 1'd0;
		12'd1269: data = 1'd0;
		12'd1270: data = 1'd0;
		12'd1271: data = 1'd0;
		12'd1272: data = 1'd0;
		12'd1273: data = 1'd0;
		12'd1274: data = 1'd1;
		12'd1275: data = 1'd1;
		12'd1276: data = 1'd0;
		12'd1277: data = 1'd1;
		12'd1278: data = 1'd0;
		12'd1279: data = 1'd1;
		12'd1280: data = 1'd0;
		12'd1281: data = 1'd0;
		12'd1282: data = 1'd0;
		12'd1283: data = 1'd1;
		12'd1284: data = 1'd0;
		12'd1285: data = 1'd1;
		12'd1286: data = 1'd0;
		12'd1287: data = 1'd1;
		12'd1288: data = 1'd1;
		12'd1289: data = 1'd0;
		12'd1290: data = 1'd1;
		12'd1291: data = 1'd0;
		12'd1292: data = 1'd0;
		12'd1293: data = 1'd1;
		12'd1294: data = 1'd0;
		12'd1295: data = 1'd0;
		12'd1296: data = 1'd1;
		12'd1297: data = 1'd1;
		12'd1298: data = 1'd0;
		12'd1299: data = 1'd1;
		12'd1300: data = 1'd0;
		12'd1301: data = 1'd1;
		12'd1302: data = 1'd0;
		12'd1303: data = 1'd1;
		12'd1304: data = 1'd0;
		12'd1305: data = 1'd0;
		12'd1306: data = 1'd1;
		12'd1307: data = 1'd0;
		12'd1308: data = 1'd0;
		12'd1309: data = 1'd1;
		12'd1310: data = 1'd0;
		12'd1311: data = 1'd0;
		12'd1312: data = 1'd1;
		12'd1313: data = 1'd0;
		12'd1314: data = 1'd1;
		12'd1315: data = 1'd0;
		12'd1316: data = 1'd1;
		12'd1317: data = 1'd0;
		12'd1318: data = 1'd0;
		12'd1319: data = 1'd1;
		12'd1320: data = 1'd0;
		12'd1321: data = 1'd1;
		12'd1322: data = 1'd1;
		12'd1323: data = 1'd0;
		12'd1324: data = 1'd0;
		12'd1325: data = 1'd1;
		12'd1326: data = 1'd1;
		12'd1327: data = 1'd0;
		12'd1328: data = 1'd1;
		12'd1329: data = 1'd0;
		12'd1330: data = 1'd1;
		12'd1331: data = 1'd0;
		12'd1332: data = 1'd1;
		12'd1333: data = 1'd0;
		12'd1334: data = 1'd0;
		12'd1335: data = 1'd1;
		12'd1336: data = 1'd1;
		12'd1337: data = 1'd0;
		12'd1338: data = 1'd1;
		12'd1339: data = 1'd1;
		12'd1340: data = 1'd0;
		12'd1341: data = 1'd0;
		12'd1342: data = 1'd1;
		12'd1343: data = 1'd1;
		12'd1344: data = 1'd1;
		12'd1345: data = 1'd0;
		12'd1346: data = 1'd0;
		12'd1347: data = 1'd1;
		12'd1348: data = 1'd0;
		12'd1349: data = 1'd1;
		12'd1350: data = 1'd0;
		12'd1351: data = 1'd0;
		12'd1352: data = 1'd1;
		12'd1353: data = 1'd1;
		12'd1354: data = 1'd0;
		12'd1355: data = 1'd0;
		12'd1356: data = 1'd1;
		12'd1357: data = 1'd1;
		12'd1358: data = 1'd0;
		12'd1359: data = 1'd1;
		12'd1360: data = 1'd1;
		12'd1361: data = 1'd0;
		12'd1362: data = 1'd0;
		12'd1363: data = 1'd0;
		12'd1364: data = 1'd1;
		12'd1365: data = 1'd0;
		12'd1366: data = 1'd1;
		12'd1367: data = 1'd0;
		12'd1368: data = 1'd0;
		12'd1369: data = 1'd1;
		12'd1370: data = 1'd1;
		12'd1371: data = 1'd0;
		12'd1372: data = 1'd0;
		12'd1373: data = 1'd1;
		12'd1374: data = 1'd1;
		12'd1375: data = 1'd0;
		12'd1376: data = 1'd1;
		12'd1377: data = 1'd0;
		12'd1378: data = 1'd0;
		12'd1379: data = 1'd0;
		12'd1380: data = 1'd1;
		12'd1381: data = 1'd0;
		12'd1382: data = 1'd0;
		12'd1383: data = 1'd1;
		12'd1384: data = 1'd0;
		12'd1385: data = 1'd0;
		12'd1386: data = 1'd1;
		12'd1387: data = 1'd1;
		12'd1388: data = 1'd0;
		12'd1389: data = 1'd0;
		12'd1390: data = 1'd1;
		12'd1391: data = 1'd1;
		12'd1392: data = 1'd1;
		12'd1393: data = 1'd0;
		12'd1394: data = 1'd0;
		12'd1395: data = 1'd0;
		12'd1396: data = 1'd1;
		12'd1397: data = 1'd0;
		12'd1398: data = 1'd0;
		12'd1399: data = 1'd1;
		12'd1400: data = 1'd0;
		12'd1401: data = 1'd0;
		12'd1402: data = 1'd0;
		12'd1403: data = 1'd1;
		12'd1404: data = 1'd1;
		12'd1405: data = 1'd0;
		12'd1406: data = 1'd0;
		12'd1407: data = 1'd1;
		12'd1408: data = 1'd0;
		12'd1409: data = 1'd1;
		12'd1410: data = 1'd1;
		12'd1411: data = 1'd1;
		12'd1412: data = 1'd1;
		12'd1413: data = 1'd0;
		12'd1414: data = 1'd0;
		12'd1415: data = 1'd1;
		12'd1416: data = 1'd0;
		12'd1417: data = 1'd0;
		12'd1418: data = 1'd0;
		12'd1419: data = 1'd1;
		12'd1420: data = 1'd1;
		12'd1421: data = 1'd1;
		12'd1422: data = 1'd0;
		12'd1423: data = 1'd0;
		12'd1424: data = 1'd1;
		12'd1425: data = 1'd0;
		12'd1426: data = 1'd1;
		12'd1427: data = 1'd1;
		12'd1428: data = 1'd1;
		12'd1429: data = 1'd0;
		12'd1430: data = 1'd0;
		12'd1431: data = 1'd1;
		12'd1432: data = 1'd0;
		12'd1433: data = 1'd0;
		12'd1434: data = 1'd1;
		12'd1435: data = 1'd1;
		12'd1436: data = 1'd1;
		12'd1437: data = 1'd0;
		12'd1438: data = 1'd0;
		12'd1439: data = 1'd0;
		12'd1440: data = 1'd0;
		12'd1441: data = 1'd0;
		12'd1442: data = 1'd0;
		12'd1443: data = 1'd0;
		12'd1444: data = 1'd0;
		12'd1445: data = 1'd1;
		12'd1446: data = 1'd0;
		12'd1447: data = 1'd1;
		12'd1448: data = 1'd0;
		12'd1449: data = 1'd0;
		12'd1450: data = 1'd1;
		12'd1451: data = 1'd1;
		12'd1452: data = 1'd0;
		12'd1453: data = 1'd0;
		12'd1454: data = 1'd0;
		12'd1455: data = 1'd1;
		12'd1456: data = 1'd0;
		12'd1457: data = 1'd0;
		12'd1458: data = 1'd0;
		12'd1459: data = 1'd0;
		12'd1460: data = 1'd0;
		12'd1461: data = 1'd0;
		12'd1462: data = 1'd1;
		12'd1463: data = 1'd0;
		12'd1464: data = 1'd1;
		12'd1465: data = 1'd0;
		12'd1466: data = 1'd1;
		12'd1467: data = 1'd0;
		12'd1468: data = 1'd0;
		12'd1469: data = 1'd1;
		12'd1470: data = 1'd1;
		12'd1471: data = 1'd1;
		12'd1472: data = 1'd0;
		12'd1473: data = 1'd0;
		12'd1474: data = 1'd0;
		12'd1475: data = 1'd0;
		12'd1476: data = 1'd0;
		12'd1477: data = 1'd0;
		12'd1478: data = 1'd0;
		12'd1479: data = 1'd1;
		12'd1480: data = 1'd1;
		12'd1481: data = 1'd0;
		12'd1482: data = 1'd1;
		12'd1483: data = 1'd0;
		12'd1484: data = 1'd0;
		12'd1485: data = 1'd1;
		12'd1486: data = 1'd0;
		12'd1487: data = 1'd0;
		12'd1488: data = 1'd0;
		12'd1489: data = 1'd0;
		12'd1490: data = 1'd0;
		12'd1491: data = 1'd0;
		12'd1492: data = 1'd0;
		12'd1493: data = 1'd0;
		12'd1494: data = 1'd0;
		12'd1495: data = 1'd0;
		12'd1496: data = 1'd0;
		12'd1497: data = 1'd1;
		12'd1498: data = 1'd0;
		12'd1499: data = 1'd1;
		12'd1500: data = 1'd0;
		12'd1501: data = 1'd1;
		12'd1502: data = 1'd0;
		12'd1503: data = 1'd0;
		12'd1504: data = 1'd0;
		12'd1505: data = 1'd0;
		12'd1506: data = 1'd0;
		12'd1507: data = 1'd0;
		12'd1508: data = 1'd0;
		12'd1509: data = 1'd0;
		12'd1510: data = 1'd0;
		12'd1511: data = 1'd0;
		12'd1512: data = 1'd0;
		12'd1513: data = 1'd0;
		12'd1514: data = 1'd1;
		12'd1515: data = 1'd0;
		12'd1516: data = 1'd1;
		12'd1517: data = 1'd1;
		12'd1518: data = 1'd1;
		12'd1519: data = 1'd0;
		12'd1520: data = 1'd0;
		12'd1521: data = 1'd0;
		12'd1522: data = 1'd0;
		12'd1523: data = 1'd0;
		12'd1524: data = 1'd0;
		12'd1525: data = 1'd0;
		12'd1526: data = 1'd0;
		12'd1527: data = 1'd0;
		12'd1528: data = 1'd0;
		12'd1529: data = 1'd0;
		12'd1530: data = 1'd1;
		12'd1531: data = 1'd0;
		12'd1532: data = 1'd1;
		12'd1533: data = 1'd0;
		12'd1534: data = 1'd1;
		12'd1535: data = 1'd0;
		12'd1536: data = 1'd0;
		12'd1537: data = 1'd0;
		12'd1538: data = 1'd0;
		12'd1539: data = 1'd0;
		12'd1540: data = 1'd0;
		12'd1541: data = 1'd0;
		12'd1542: data = 1'd0;
		12'd1543: data = 1'd0;
		12'd1544: data = 1'd1;
		12'd1545: data = 1'd1;
		12'd1546: data = 1'd0;
		12'd1547: data = 1'd1;
		12'd1548: data = 1'd1;
		12'd1549: data = 1'd0;
		12'd1550: data = 1'd0;
		12'd1551: data = 1'd0;
		12'd1552: data = 1'd0;
		12'd1553: data = 1'd0;
		12'd1554: data = 1'd0;
		12'd1555: data = 1'd0;
		12'd1556: data = 1'd0;
		12'd1557: data = 1'd0;
		12'd1558: data = 1'd0;
		12'd1559: data = 1'd0;
		12'd1560: data = 1'd1;
		12'd1561: data = 1'd1;
		12'd1562: data = 1'd0;
		12'd1563: data = 1'd1;
		12'd1564: data = 1'd0;
		12'd1565: data = 1'd0;
		12'd1566: data = 1'd1;
		12'd1567: data = 1'd1;
		12'd1568: data = 1'd0;
		12'd1569: data = 1'd0;
		12'd1570: data = 1'd0;
		12'd1571: data = 1'd0;
		12'd1572: data = 1'd0;
		12'd1573: data = 1'd0;
		12'd1574: data = 1'd0;
		12'd1575: data = 1'd0;
		12'd1576: data = 1'd1;
		12'd1577: data = 1'd0;
		12'd1578: data = 1'd0;
		12'd1579: data = 1'd1;
		12'd1580: data = 1'd0;
		12'd1581: data = 1'd0;
		12'd1582: data = 1'd1;
		12'd1583: data = 1'd0;
		12'd1584: data = 1'd0;
		12'd1585: data = 1'd0;
		12'd1586: data = 1'd0;
		12'd1587: data = 1'd0;
		12'd1588: data = 1'd0;
		12'd1589: data = 1'd0;
		12'd1590: data = 1'd0;
		12'd1591: data = 1'd0;
		12'd1592: data = 1'd1;
		12'd1593: data = 1'd0;
		12'd1594: data = 1'd1;
		12'd1595: data = 1'd1;
		12'd1596: data = 1'd0;
		12'd1597: data = 1'd0;
		12'd1598: data = 1'd1;
		12'd1599: data = 1'd1;
		12'd1600: data = 1'd0;
		12'd1601: data = 1'd0;
		12'd1602: data = 1'd0;
		12'd1603: data = 1'd0;
		12'd1604: data = 1'd0;
		12'd1605: data = 1'd0;
		12'd1606: data = 1'd0;
		12'd1607: data = 1'd0;
		12'd1608: data = 1'd1;
		12'd1609: data = 1'd1;
		12'd1610: data = 1'd0;
		12'd1611: data = 1'd0;
		12'd1612: data = 1'd1;
		12'd1613: data = 1'd0;
		12'd1614: data = 1'd0;
		12'd1615: data = 1'd0;
		12'd1616: data = 1'd0;
		12'd1617: data = 1'd0;
		12'd1618: data = 1'd0;
		12'd1619: data = 1'd0;
		12'd1620: data = 1'd0;
		12'd1621: data = 1'd0;
		12'd1622: data = 1'd0;
		12'd1623: data = 1'd0;
		12'd1624: data = 1'd0;
		12'd1625: data = 1'd1;
		12'd1626: data = 1'd1;
		12'd1627: data = 1'd0;
		12'd1628: data = 1'd0;
		12'd1629: data = 1'd1;
		12'd1630: data = 1'd1;
		12'd1631: data = 1'd0;
		12'd1632: data = 1'd0;
		12'd1633: data = 1'd0;
		12'd1634: data = 1'd0;
		12'd1635: data = 1'd0;
		12'd1636: data = 1'd0;
		12'd1637: data = 1'd0;
		12'd1638: data = 1'd0;
		12'd1639: data = 1'd0;
		12'd1640: data = 1'd0;
		12'd1641: data = 1'd0;
		12'd1642: data = 1'd1;
		12'd1643: data = 1'd1;
		12'd1644: data = 1'd0;
		12'd1645: data = 1'd0;
		12'd1646: data = 1'd1;
		12'd1647: data = 1'd1;
		12'd1648: data = 1'd0;
		12'd1649: data = 1'd0;
		12'd1650: data = 1'd0;
		12'd1651: data = 1'd0;
		12'd1652: data = 1'd0;
		12'd1653: data = 1'd0;
		12'd1654: data = 1'd0;
		12'd1655: data = 1'd0;
		12'd1656: data = 1'd0;
		12'd1657: data = 1'd0;
		12'd1658: data = 1'd0;
		12'd1659: data = 1'd1;
		12'd1660: data = 1'd1;
		12'd1661: data = 1'd0;
		12'd1662: data = 1'd0;
		12'd1663: data = 1'd1;
		12'd1664: data = 1'd0;
		12'd1665: data = 1'd0;
		12'd1666: data = 1'd0;
		12'd1667: data = 1'd0;
		12'd1668: data = 1'd0;
		12'd1669: data = 1'd0;
		12'd1670: data = 1'd0;
		12'd1671: data = 1'd0;
		12'd1672: data = 1'd0;
		12'd1673: data = 1'd0;
		12'd1674: data = 1'd0;
		12'd1675: data = 1'd0;
		12'd1676: data = 1'd1;
		12'd1677: data = 1'd1;
		12'd1678: data = 1'd0;
		12'd1679: data = 1'd1;
		12'd1680: data = 1'd0;
		12'd1681: data = 1'd0;
		12'd1682: data = 1'd0;
		12'd1683: data = 1'd0;
		12'd1684: data = 1'd0;
		12'd1685: data = 1'd0;
		12'd1686: data = 1'd0;
		12'd1687: data = 1'd0;
		12'd1688: data = 1'd0;
		12'd1689: data = 1'd0;
		12'd1690: data = 1'd0;
		12'd1691: data = 1'd0;
		12'd1692: data = 1'd1;
		12'd1693: data = 1'd1;
		12'd1694: data = 1'd1;
		12'd1695: data = 1'd0;
		12'd1696: data = 1'd0;
		12'd1697: data = 1'd0;
		12'd1698: data = 1'd0;
		12'd1699: data = 1'd0;
		12'd1700: data = 1'd0;
		12'd1701: data = 1'd0;
		12'd1702: data = 1'd0;
		12'd1703: data = 1'd0;
		12'd1704: data = 1'd0;
		12'd1705: data = 1'd0;
		12'd1706: data = 1'd0;
		12'd1707: data = 1'd1;
		12'd1708: data = 1'd1;
		12'd1709: data = 1'd1;
		12'd1710: data = 1'd0;
		12'd1711: data = 1'd0;
		12'd1712: data = 1'd0;
		12'd1713: data = 1'd0;
		12'd1714: data = 1'd0;
		12'd1715: data = 1'd0;
		12'd1716: data = 1'd0;
		12'd1717: data = 1'd0;
		12'd1718: data = 1'd0;
		12'd1719: data = 1'd0;
		12'd1720: data = 1'd0;
		12'd1721: data = 1'd0;
		12'd1722: data = 1'd0;
		12'd1723: data = 1'd1;
		12'd1724: data = 1'd1;
		12'd1725: data = 1'd0;
		12'd1726: data = 1'd0;
		12'd1727: data = 1'd1;
		12'd1728: data = 1'd0;
		12'd1729: data = 1'd0;
		12'd1730: data = 1'd0;
		12'd1731: data = 1'd0;
		12'd1732: data = 1'd0;
		12'd1733: data = 1'd0;
		12'd1734: data = 1'd0;
		12'd1735: data = 1'd0;
		12'd1736: data = 1'd0;
		12'd1737: data = 1'd0;
		12'd1738: data = 1'd0;
		12'd1739: data = 1'd1;
		12'd1740: data = 1'd0;
		12'd1741: data = 1'd0;
		12'd1742: data = 1'd1;
		12'd1743: data = 1'd0;
		12'd1744: data = 1'd0;
		12'd1745: data = 1'd0;
		12'd1746: data = 1'd0;
		12'd1747: data = 1'd0;
		12'd1748: data = 1'd0;
		12'd1749: data = 1'd0;
		12'd1750: data = 1'd0;
		12'd1751: data = 1'd0;
		12'd1752: data = 1'd0;
		12'd1753: data = 1'd0;
		12'd1754: data = 1'd0;
		12'd1755: data = 1'd1;
		12'd1756: data = 1'd0;
		12'd1757: data = 1'd1;
		12'd1758: data = 1'd0;
		12'd1759: data = 1'd1;
		12'd1760: data = 1'd0;
		12'd1761: data = 1'd0;
		12'd1762: data = 1'd0;
		12'd1763: data = 1'd0;
		12'd1764: data = 1'd0;
		12'd1765: data = 1'd0;
		12'd1766: data = 1'd0;
		12'd1767: data = 1'd0;
		12'd1768: data = 1'd0;
		12'd1769: data = 1'd0;
		12'd1770: data = 1'd0;
		12'd1771: data = 1'd1;
		12'd1772: data = 1'd0;
		12'd1773: data = 1'd1;
		12'd1774: data = 1'd0;
		12'd1775: data = 1'd1;
		12'd1776: data = 1'd0;
		12'd1777: data = 1'd0;
		12'd1778: data = 1'd0;
		12'd1779: data = 1'd0;
		12'd1780: data = 1'd0;
		12'd1781: data = 1'd0;
		12'd1782: data = 1'd0;
		12'd1783: data = 1'd0;
		12'd1784: data = 1'd0;
		12'd1785: data = 1'd0;
		12'd1786: data = 1'd0;
		12'd1787: data = 1'd1;
		12'd1788: data = 1'd0;
		12'd1789: data = 1'd1;
		12'd1790: data = 1'd1;
		12'd1791: data = 1'd0;
		12'd1792: data = 1'd0;
		12'd1793: data = 1'd0;
		12'd1794: data = 1'd0;
		12'd1795: data = 1'd0;
		12'd1796: data = 1'd0;
		12'd1797: data = 1'd0;
		12'd1798: data = 1'd0;
		12'd1799: data = 1'd0;
		12'd1800: data = 1'd0;
		12'd1801: data = 1'd0;
		12'd1802: data = 1'd0;
		12'd1803: data = 1'd0;
		12'd1804: data = 1'd0;
		12'd1805: data = 1'd0;
		12'd1806: data = 1'd0;
		12'd1807: data = 1'd0;
		12'd1808: data = 1'd0;
		12'd1809: data = 1'd0;
		12'd1810: data = 1'd0;
		12'd1811: data = 1'd0;
		12'd1812: data = 1'd0;
		12'd1813: data = 1'd0;
		12'd1814: data = 1'd0;
		12'd1815: data = 1'd0;
		12'd1816: data = 1'd0;
		12'd1817: data = 1'd0;
		12'd1818: data = 1'd0;
		12'd1819: data = 1'd0;
		12'd1820: data = 1'd0;
		12'd1821: data = 1'd0;
		12'd1822: data = 1'd0;
		12'd1823: data = 1'd1;
		12'd1824: data = 1'd0;
		12'd1825: data = 1'd0;
		12'd1826: data = 1'd0;
		12'd1827: data = 1'd0;
		12'd1828: data = 1'd0;
		12'd1829: data = 1'd0;
		12'd1830: data = 1'd0;
		12'd1831: data = 1'd0;
		12'd1832: data = 1'd0;
		12'd1833: data = 1'd0;
		12'd1834: data = 1'd0;
		12'd1835: data = 1'd0;
		12'd1836: data = 1'd0;
		12'd1837: data = 1'd0;
		12'd1838: data = 1'd1;
		12'd1839: data = 1'd0;
		12'd1840: data = 1'd0;
		12'd1841: data = 1'd0;
		12'd1842: data = 1'd0;
		12'd1843: data = 1'd0;
		12'd1844: data = 1'd0;
		12'd1845: data = 1'd0;
		12'd1846: data = 1'd0;
		12'd1847: data = 1'd0;
		12'd1848: data = 1'd0;
		12'd1849: data = 1'd0;
		12'd1850: data = 1'd0;
		12'd1851: data = 1'd0;
		12'd1852: data = 1'd0;
		12'd1853: data = 1'd1;
		12'd1854: data = 1'd0;
		12'd1855: data = 1'd1;
		12'd1856: data = 1'd0;
		12'd1857: data = 1'd0;
		12'd1858: data = 1'd0;
		12'd1859: data = 1'd0;
		12'd1860: data = 1'd0;
		12'd1861: data = 1'd0;
		12'd1862: data = 1'd0;
		12'd1863: data = 1'd0;
		12'd1864: data = 1'd0;
		12'd1865: data = 1'd0;
		12'd1866: data = 1'd0;
		12'd1867: data = 1'd0;
		12'd1868: data = 1'd0;
		12'd1869: data = 1'd1;
		12'd1870: data = 1'd0;
		12'd1871: data = 1'd1;
		12'd1872: data = 1'd0;
		12'd1873: data = 1'd0;
		12'd1874: data = 1'd0;
		12'd1875: data = 1'd0;
		12'd1876: data = 1'd0;
		12'd1877: data = 1'd0;
		12'd1878: data = 1'd0;
		12'd1879: data = 1'd0;
		12'd1880: data = 1'd0;
		12'd1881: data = 1'd0;
		12'd1882: data = 1'd0;
		12'd1883: data = 1'd0;
		12'd1884: data = 1'd0;
		12'd1885: data = 1'd1;
		12'd1886: data = 1'd0;
		12'd1887: data = 1'd1;
		12'd1888: data = 1'd0;
		12'd1889: data = 1'd0;
		12'd1890: data = 1'd0;
		12'd1891: data = 1'd0;
		12'd1892: data = 1'd0;
		12'd1893: data = 1'd0;
		12'd1894: data = 1'd0;
		12'd1895: data = 1'd0;
		12'd1896: data = 1'd0;
		12'd1897: data = 1'd0;
		12'd1898: data = 1'd0;
		12'd1899: data = 1'd0;
		12'd1900: data = 1'd0;
		12'd1901: data = 1'd1;
		12'd1902: data = 1'd0;
		12'd1903: data = 1'd0;
		12'd1904: data = 1'd0;
		12'd1905: data = 1'd0;
		12'd1906: data = 1'd0;
		12'd1907: data = 1'd0;
		12'd1908: data = 1'd0;
		12'd1909: data = 1'd0;
		12'd1910: data = 1'd0;
		12'd1911: data = 1'd0;
		12'd1912: data = 1'd0;
		12'd1913: data = 1'd0;
		12'd1914: data = 1'd0;
		12'd1915: data = 1'd0;
		12'd1916: data = 1'd0;
		12'd1917: data = 1'd0;
		12'd1918: data = 1'd1;
		12'd1919: data = 1'd0;
		12'd1920: data = 1'd0;
		12'd1921: data = 1'd0;
		12'd1922: data = 1'd0;
		12'd1923: data = 1'd0;
		12'd1924: data = 1'd0;
		12'd1925: data = 1'd0;
		12'd1926: data = 1'd0;
		12'd1927: data = 1'd0;
		12'd1928: data = 1'd0;
		12'd1929: data = 1'd0;
		12'd1930: data = 1'd0;
		12'd1931: data = 1'd0;
		12'd1932: data = 1'd0;
		12'd1933: data = 1'd0;
		12'd1934: data = 1'd1;
		12'd1935: data = 1'd0;
		12'd1936: data = 1'd0;
		12'd1937: data = 1'd0;
		12'd1938: data = 1'd0;
		12'd1939: data = 1'd0;
		12'd1940: data = 1'd0;
		12'd1941: data = 1'd0;
		12'd1942: data = 1'd0;
		12'd1943: data = 1'd0;
		12'd1944: data = 1'd0;
		12'd1945: data = 1'd0;
		12'd1946: data = 1'd0;
		12'd1947: data = 1'd0;
		12'd1948: data = 1'd0;
		12'd1949: data = 1'd0;
		12'd1950: data = 1'd0;
		12'd1951: data = 1'd1;
		12'd1952: data = 1'd0;
		12'd1953: data = 1'd0;
		12'd1954: data = 1'd0;
		12'd1955: data = 1'd0;
		12'd1956: data = 1'd0;
		12'd1957: data = 1'd0;
		12'd1958: data = 1'd0;
		12'd1959: data = 1'd0;
		12'd1960: data = 1'd0;
		12'd1961: data = 1'd0;
		12'd1962: data = 1'd0;
		12'd1963: data = 1'd0;
		12'd1964: data = 1'd0;
		12'd1965: data = 1'd0;
		12'd1966: data = 1'd0;
		12'd1967: data = 1'd1;
		12'd1968: data = 1'd0;
		12'd1969: data = 1'd0;
		12'd1970: data = 1'd0;
		12'd1971: data = 1'd0;
		12'd1972: data = 1'd0;
		12'd1973: data = 1'd0;
		12'd1974: data = 1'd0;
		12'd1975: data = 1'd0;
		12'd1976: data = 1'd0;
		12'd1977: data = 1'd0;
		12'd1978: data = 1'd0;
		12'd1979: data = 1'd0;
		12'd1980: data = 1'd0;
		12'd1981: data = 1'd0;
		12'd1982: data = 1'd1;
		12'd1983: data = 1'd0;
		12'd1984: data = 1'd0;
		12'd1985: data = 1'd0;
		12'd1986: data = 1'd0;
		12'd1987: data = 1'd0;
		12'd1988: data = 1'd0;
		12'd1989: data = 1'd0;
		12'd1990: data = 1'd0;
		12'd1991: data = 1'd0;
		12'd1992: data = 1'd0;
		12'd1993: data = 1'd0;
		12'd1994: data = 1'd0;
		12'd1995: data = 1'd0;
		12'd1996: data = 1'd1;
		12'd1997: data = 1'd1;
		12'd1998: data = 1'd0;
		12'd1999: data = 1'd0;
		12'd2000: data = 1'd0;
		12'd2001: data = 1'd0;
		12'd2002: data = 1'd0;
		12'd2003: data = 1'd0;
		12'd2004: data = 1'd0;
		12'd2005: data = 1'd0;
		12'd2006: data = 1'd0;
		12'd2007: data = 1'd0;
		12'd2008: data = 1'd0;
		12'd2009: data = 1'd0;
		12'd2010: data = 1'd0;
		12'd2011: data = 1'd1;
		12'd2012: data = 1'd0;
		12'd2013: data = 1'd1;
		12'd2014: data = 1'd1;
		12'd2015: data = 1'd0;
		12'd2016: data = 1'd0;
		12'd2017: data = 1'd0;
		12'd2018: data = 1'd0;
		12'd2019: data = 1'd0;
		12'd2020: data = 1'd0;
		12'd2021: data = 1'd0;
		12'd2022: data = 1'd0;
		12'd2023: data = 1'd0;
		12'd2024: data = 1'd0;
		12'd2025: data = 1'd0;
		12'd2026: data = 1'd0;
		12'd2027: data = 1'd1;
		12'd2028: data = 1'd0;
		12'd2029: data = 1'd1;
		12'd2030: data = 1'd0;
		12'd2031: data = 1'd1;
		12'd2032: data = 1'd0;
		12'd2033: data = 1'd0;
		12'd2034: data = 1'd0;
		12'd2035: data = 1'd0;
		12'd2036: data = 1'd0;
		12'd2037: data = 1'd0;
		12'd2038: data = 1'd0;
		12'd2039: data = 1'd0;
		12'd2040: data = 1'd0;
		12'd2041: data = 1'd0;
		12'd2042: data = 1'd0;
		12'd2043: data = 1'd1;
		12'd2044: data = 1'd0;
		12'd2045: data = 1'd1;
		12'd2046: data = 1'd0;
		12'd2047: data = 1'd1;
		12'd2048: data = 1'd0;
		12'd2049: data = 1'd0;
		12'd2050: data = 1'd0;
		12'd2051: data = 1'd0;
		12'd2052: data = 1'd0;
		12'd2053: data = 1'd0;
		12'd2054: data = 1'd0;
		12'd2055: data = 1'd0;
		12'd2056: data = 1'd0;
		12'd2057: data = 1'd0;
		12'd2058: data = 1'd0;
		12'd2059: data = 1'd0;
		12'd2060: data = 1'd0;
		12'd2061: data = 1'd0;
		12'd2062: data = 1'd0;
		12'd2063: data = 1'd0;
		12'd2064: data = 1'd0;
		12'd2065: data = 1'd0;
		12'd2066: data = 1'd0;
		12'd2067: data = 1'd0;
		12'd2068: data = 1'd0;
		12'd2069: data = 1'd0;
		12'd2070: data = 1'd0;
		12'd2071: data = 1'd0;
		12'd2072: data = 1'd0;
		12'd2073: data = 1'd0;
		12'd2074: data = 1'd0;
		12'd2075: data = 1'd0;
		12'd2076: data = 1'd0;
		12'd2077: data = 1'd0;
		12'd2078: data = 1'd0;
		12'd2079: data = 1'd0;
		12'd2080: data = 1'd0;
		12'd2081: data = 1'd0;
		12'd2082: data = 1'd0;
		12'd2083: data = 1'd0;
		12'd2084: data = 1'd0;
		12'd2085: data = 1'd0;
		12'd2086: data = 1'd0;
		12'd2087: data = 1'd0;
		12'd2088: data = 1'd0;
		12'd2089: data = 1'd0;
		12'd2090: data = 1'd0;
		12'd2091: data = 1'd0;
		12'd2092: data = 1'd0;
		12'd2093: data = 1'd0;
		12'd2094: data = 1'd0;
		12'd2095: data = 1'd1;
		12'd2096: data = 1'd0;
		12'd2097: data = 1'd0;
		12'd2098: data = 1'd0;
		12'd2099: data = 1'd0;
		12'd2100: data = 1'd0;
		12'd2101: data = 1'd0;
		12'd2102: data = 1'd0;
		12'd2103: data = 1'd0;
		12'd2104: data = 1'd0;
		12'd2105: data = 1'd0;
		12'd2106: data = 1'd0;
		12'd2107: data = 1'd0;
		12'd2108: data = 1'd0;
		12'd2109: data = 1'd0;
		12'd2110: data = 1'd1;
		12'd2111: data = 1'd0;
		12'd2112: data = 1'd0;
		12'd2113: data = 1'd0;
		12'd2114: data = 1'd0;
		12'd2115: data = 1'd0;
		12'd2116: data = 1'd0;
		12'd2117: data = 1'd0;
		12'd2118: data = 1'd0;
		12'd2119: data = 1'd0;
		12'd2120: data = 1'd0;
		12'd2121: data = 1'd0;
		12'd2122: data = 1'd0;
		12'd2123: data = 1'd0;
		12'd2124: data = 1'd0;
		12'd2125: data = 1'd1;
		12'd2126: data = 1'd0;
		12'd2127: data = 1'd1;
		12'd2128: data = 1'd0;
		12'd2129: data = 1'd0;
		12'd2130: data = 1'd0;
		12'd2131: data = 1'd0;
		12'd2132: data = 1'd0;
		12'd2133: data = 1'd0;
		12'd2134: data = 1'd0;
		12'd2135: data = 1'd0;
		12'd2136: data = 1'd0;
		12'd2137: data = 1'd0;
		12'd2138: data = 1'd0;
		12'd2139: data = 1'd0;
		12'd2140: data = 1'd0;
		12'd2141: data = 1'd1;
		12'd2142: data = 1'd1;
		12'd2143: data = 1'd0;
		12'd2144: data = 1'd0;
		12'd2145: data = 1'd0;
		12'd2146: data = 1'd0;
		12'd2147: data = 1'd0;
		12'd2148: data = 1'd0;
		12'd2149: data = 1'd0;
		12'd2150: data = 1'd0;
		12'd2151: data = 1'd0;
		12'd2152: data = 1'd0;
		12'd2153: data = 1'd0;
		12'd2154: data = 1'd0;
		12'd2155: data = 1'd0;
		12'd2156: data = 1'd0;
		12'd2157: data = 1'd0;
		12'd2158: data = 1'd1;
		12'd2159: data = 1'd1;
		12'd2160: data = 1'd0;
		12'd2161: data = 1'd0;
		12'd2162: data = 1'd0;
		12'd2163: data = 1'd0;
		12'd2164: data = 1'd0;
		12'd2165: data = 1'd0;
		12'd2166: data = 1'd0;
		12'd2167: data = 1'd0;
		12'd2168: data = 1'd0;
		12'd2169: data = 1'd0;
		12'd2170: data = 1'd0;
		12'd2171: data = 1'd0;
		12'd2172: data = 1'd0;
		12'd2173: data = 1'd0;
		12'd2174: data = 1'd0;
		12'd2175: data = 1'd1;
		12'd2176: data = 1'd0;
		12'd2177: data = 1'd0;
		12'd2178: data = 1'd0;
		12'd2179: data = 1'd0;
		12'd2180: data = 1'd0;
		12'd2181: data = 1'd0;
		12'd2182: data = 1'd0;
		12'd2183: data = 1'd0;
		12'd2184: data = 1'd0;
		12'd2185: data = 1'd0;
		12'd2186: data = 1'd0;
		12'd2187: data = 1'd0;
		12'd2188: data = 1'd0;
		12'd2189: data = 1'd0;
		12'd2190: data = 1'd0;
		12'd2191: data = 1'd1;
		12'd2192: data = 1'd0;
		12'd2193: data = 1'd0;
		12'd2194: data = 1'd0;
		12'd2195: data = 1'd0;
		12'd2196: data = 1'd0;
		12'd2197: data = 1'd0;
		12'd2198: data = 1'd0;
		12'd2199: data = 1'd0;
		12'd2200: data = 1'd0;
		12'd2201: data = 1'd0;
		12'd2202: data = 1'd0;
		12'd2203: data = 1'd0;
		12'd2204: data = 1'd0;
		12'd2205: data = 1'd0;
		12'd2206: data = 1'd0;
		12'd2207: data = 1'd0;
		12'd2208: data = 1'd0;
		12'd2209: data = 1'd0;
		12'd2210: data = 1'd0;
		12'd2211: data = 1'd0;
		12'd2212: data = 1'd0;
		12'd2213: data = 1'd0;
		12'd2214: data = 1'd0;
		12'd2215: data = 1'd0;
		12'd2216: data = 1'd0;
		12'd2217: data = 1'd0;
		12'd2218: data = 1'd0;
		12'd2219: data = 1'd0;
		12'd2220: data = 1'd0;
		12'd2221: data = 1'd0;
		12'd2222: data = 1'd0;
		12'd2223: data = 1'd0;
		12'd2224: data = 1'd0;
		12'd2225: data = 1'd0;
		12'd2226: data = 1'd0;
		12'd2227: data = 1'd0;
		12'd2228: data = 1'd0;
		12'd2229: data = 1'd0;
		12'd2230: data = 1'd0;
		12'd2231: data = 1'd0;
		12'd2232: data = 1'd0;
		12'd2233: data = 1'd0;
		12'd2234: data = 1'd0;
		12'd2235: data = 1'd0;
		12'd2236: data = 1'd0;
		12'd2237: data = 1'd0;
		12'd2238: data = 1'd0;
		12'd2239: data = 1'd1;
		12'd2240: data = 1'd0;
		12'd2241: data = 1'd0;
		12'd2242: data = 1'd0;
		12'd2243: data = 1'd0;
		12'd2244: data = 1'd0;
		12'd2245: data = 1'd0;
		12'd2246: data = 1'd0;
		12'd2247: data = 1'd0;
		12'd2248: data = 1'd0;
		12'd2249: data = 1'd0;
		12'd2250: data = 1'd0;
		12'd2251: data = 1'd0;
		12'd2252: data = 1'd1;
		12'd2253: data = 1'd1;
		12'd2254: data = 1'd0;
		12'd2255: data = 1'd0;
		12'd2256: data = 1'd0;
		12'd2257: data = 1'd0;
		12'd2258: data = 1'd0;
		12'd2259: data = 1'd0;
		12'd2260: data = 1'd0;
		12'd2261: data = 1'd0;
		12'd2262: data = 1'd0;
		12'd2263: data = 1'd0;
		12'd2264: data = 1'd0;
		12'd2265: data = 1'd0;
		12'd2266: data = 1'd0;
		12'd2267: data = 1'd0;
		12'd2268: data = 1'd0;
		12'd2269: data = 1'd1;
		12'd2270: data = 1'd1;
		12'd2271: data = 1'd0;
		12'd2272: data = 1'd0;
		12'd2273: data = 1'd0;
		12'd2274: data = 1'd0;
		12'd2275: data = 1'd0;
		12'd2276: data = 1'd0;
		12'd2277: data = 1'd0;
		12'd2278: data = 1'd0;
		12'd2279: data = 1'd0;
		12'd2280: data = 1'd0;
		12'd2281: data = 1'd0;
		12'd2282: data = 1'd0;
		12'd2283: data = 1'd0;
		12'd2284: data = 1'd1;
		12'd2285: data = 1'd0;
		12'd2286: data = 1'd1;
		12'd2287: data = 1'd1;
		12'd2288: data = 1'd0;
		12'd2289: data = 1'd0;
		12'd2290: data = 1'd0;
		12'd2291: data = 1'd0;
		12'd2292: data = 1'd0;
		12'd2293: data = 1'd0;
		12'd2294: data = 1'd0;
		12'd2295: data = 1'd0;
		12'd2296: data = 1'd0;
		12'd2297: data = 1'd0;
		12'd2298: data = 1'd0;
		12'd2299: data = 1'd0;
		12'd2300: data = 1'd1;
		12'd2301: data = 1'd0;
		12'd2302: data = 1'd1;
		12'd2303: data = 1'd0;
		12'd2304: data = 1'd0;
		12'd2305: data = 1'd0;
		12'd2306: data = 1'd0;
		12'd2307: data = 1'd0;
		12'd2308: data = 1'd0;
		12'd2309: data = 1'd0;
		12'd2310: data = 1'd0;
		12'd2311: data = 1'd0;
		12'd2312: data = 1'd0;
		12'd2313: data = 1'd0;
		12'd2314: data = 1'd0;
		12'd2315: data = 1'd0;
		12'd2316: data = 1'd0;
		12'd2317: data = 1'd0;
		12'd2318: data = 1'd0;
		12'd2319: data = 1'd0;
		12'd2320: data = 1'd0;
		12'd2321: data = 1'd0;
		12'd2322: data = 1'd0;
		12'd2323: data = 1'd0;
		12'd2324: data = 1'd0;
		12'd2325: data = 1'd0;
		12'd2326: data = 1'd0;
		12'd2327: data = 1'd0;
		12'd2328: data = 1'd0;
		12'd2329: data = 1'd0;
		12'd2330: data = 1'd0;
		12'd2331: data = 1'd0;
		12'd2332: data = 1'd0;
		12'd2333: data = 1'd0;
		12'd2334: data = 1'd0;
		12'd2335: data = 1'd1;
		12'd2336: data = 1'd0;
		12'd2337: data = 1'd0;
		12'd2338: data = 1'd0;
		12'd2339: data = 1'd0;
		12'd2340: data = 1'd0;
		12'd2341: data = 1'd0;
		12'd2342: data = 1'd0;
		12'd2343: data = 1'd0;
		12'd2344: data = 1'd0;
		12'd2345: data = 1'd0;
		12'd2346: data = 1'd0;
		12'd2347: data = 1'd0;
		12'd2348: data = 1'd0;
		12'd2349: data = 1'd0;
		12'd2350: data = 1'd1;
		12'd2351: data = 1'd0;
		12'd2352: data = 1'd0;
		12'd2353: data = 1'd0;
		12'd2354: data = 1'd0;
		12'd2355: data = 1'd0;
		12'd2356: data = 1'd0;
		12'd2357: data = 1'd0;
		12'd2358: data = 1'd0;
		12'd2359: data = 1'd0;
		12'd2360: data = 1'd0;
		12'd2361: data = 1'd0;
		12'd2362: data = 1'd0;
		12'd2363: data = 1'd0;
		12'd2364: data = 1'd0;
		12'd2365: data = 1'd1;
		12'd2366: data = 1'd0;
		12'd2367: data = 1'd0;
		12'd2368: data = 1'd0;
		12'd2369: data = 1'd0;
		12'd2370: data = 1'd0;
		12'd2371: data = 1'd0;
		12'd2372: data = 1'd0;
		12'd2373: data = 1'd0;
		12'd2374: data = 1'd0;
		12'd2375: data = 1'd0;
		12'd2376: data = 1'd0;
		12'd2377: data = 1'd0;
		12'd2378: data = 1'd0;
		12'd2379: data = 1'd0;
		12'd2380: data = 1'd0;
		12'd2381: data = 1'd1;
		12'd2382: data = 1'd0;
		12'd2383: data = 1'd1;
		12'd2384: data = 1'd0;
		12'd2385: data = 1'd0;
		12'd2386: data = 1'd0;
		12'd2387: data = 1'd0;
		12'd2388: data = 1'd0;
		12'd2389: data = 1'd0;
		12'd2390: data = 1'd0;
		12'd2391: data = 1'd0;
		12'd2392: data = 1'd0;
		12'd2393: data = 1'd0;
		12'd2394: data = 1'd1;
		12'd2395: data = 1'd0;
		12'd2396: data = 1'd1;
		12'd2397: data = 1'd0;
		12'd2398: data = 1'd1;
		12'd2399: data = 1'd1;
		12'd2400: data = 1'd0;
		12'd2401: data = 1'd0;
		12'd2402: data = 1'd0;
		12'd2403: data = 1'd0;
		12'd2404: data = 1'd0;
		12'd2405: data = 1'd0;
		12'd2406: data = 1'd1;
		12'd2407: data = 1'd0;
		12'd2408: data = 1'd1;
		12'd2409: data = 1'd1;
		12'd2410: data = 1'd0;
		12'd2411: data = 1'd1;
		12'd2412: data = 1'd1;
		12'd2413: data = 1'd0;
		12'd2414: data = 1'd0;
		12'd2415: data = 1'd0;
		12'd2416: data = 1'd0;
		12'd2417: data = 1'd0;
		12'd2418: data = 1'd0;
		12'd2419: data = 1'd0;
		12'd2420: data = 1'd1;
		12'd2421: data = 1'd1;
		12'd2422: data = 1'd1;
		12'd2423: data = 1'd1;
		12'd2424: data = 1'd1;
		12'd2425: data = 1'd0;
		12'd2426: data = 1'd1;
		12'd2427: data = 1'd1;
		12'd2428: data = 1'd0;
		12'd2429: data = 1'd1;
		12'd2430: data = 1'd1;
		12'd2431: data = 1'd0;
		12'd2432: data = 1'd0;
		12'd2433: data = 1'd0;
		12'd2434: data = 1'd0;
		12'd2435: data = 1'd0;
		12'd2436: data = 1'd0;
		12'd2437: data = 1'd1;
		12'd2438: data = 1'd0;
		12'd2439: data = 1'd1;
		12'd2440: data = 1'd0;
		12'd2441: data = 1'd1;
		12'd2442: data = 1'd0;
		12'd2443: data = 1'd0;
		12'd2444: data = 1'd1;
		12'd2445: data = 1'd1;
		12'd2446: data = 1'd0;
		12'd2447: data = 1'd1;
		12'd2448: data = 1'd0;
		12'd2449: data = 1'd0;
		12'd2450: data = 1'd0;
		12'd2451: data = 1'd0;
		12'd2452: data = 1'd0;
		12'd2453: data = 1'd0;
		12'd2454: data = 1'd0;
		12'd2455: data = 1'd1;
		12'd2456: data = 1'd0;
		12'd2457: data = 1'd0;
		12'd2458: data = 1'd1;
		12'd2459: data = 1'd1;
		12'd2460: data = 1'd0;
		12'd2461: data = 1'd0;
		12'd2462: data = 1'd1;
		12'd2463: data = 1'd0;
		12'd2464: data = 1'd0;
		12'd2465: data = 1'd0;
		12'd2466: data = 1'd0;
		12'd2467: data = 1'd0;
		12'd2468: data = 1'd0;
		12'd2469: data = 1'd1;
		12'd2470: data = 1'd1;
		12'd2471: data = 1'd1;
		12'd2472: data = 1'd0;
		12'd2473: data = 1'd0;
		12'd2474: data = 1'd1;
		12'd2475: data = 1'd0;
		12'd2476: data = 1'd1;
		12'd2477: data = 1'd1;
		12'd2478: data = 1'd0;
		12'd2479: data = 1'd1;
		12'd2480: data = 1'd0;
		12'd2481: data = 1'd0;
		12'd2482: data = 1'd0;
		12'd2483: data = 1'd0;
		12'd2484: data = 1'd0;
		12'd2485: data = 1'd0;
		12'd2486: data = 1'd1;
		12'd2487: data = 1'd1;
		12'd2488: data = 1'd0;
		12'd2489: data = 1'd1;
		12'd2490: data = 1'd1;
		12'd2491: data = 1'd0;
		12'd2492: data = 1'd0;
		12'd2493: data = 1'd1;
		12'd2494: data = 1'd1;
		12'd2495: data = 1'd1;
		12'd2496: data = 1'd0;
		12'd2497: data = 1'd0;
		12'd2498: data = 1'd0;
		12'd2499: data = 1'd0;
		12'd2500: data = 1'd0;
		12'd2501: data = 1'd0;
		12'd2502: data = 1'd0;
		12'd2503: data = 1'd0;
		12'd2504: data = 1'd0;
		12'd2505: data = 1'd1;
		12'd2506: data = 1'd0;
		12'd2507: data = 1'd0;
		12'd2508: data = 1'd0;
		12'd2509: data = 1'd0;
		12'd2510: data = 1'd1;
		12'd2511: data = 1'd1;
		12'd2512: data = 1'd0;
		12'd2513: data = 1'd0;
		12'd2514: data = 1'd0;
		12'd2515: data = 1'd0;
		12'd2516: data = 1'd0;
		12'd2517: data = 1'd0;
		12'd2518: data = 1'd1;
		12'd2519: data = 1'd1;
		12'd2520: data = 1'd0;
		12'd2521: data = 1'd0;
		12'd2522: data = 1'd0;
		12'd2523: data = 1'd1;
		12'd2524: data = 1'd0;
		12'd2525: data = 1'd0;
		12'd2526: data = 1'd0;
		12'd2527: data = 1'd0;
		12'd2528: data = 1'd0;
		12'd2529: data = 1'd0;
		12'd2530: data = 1'd0;
		12'd2531: data = 1'd0;
		12'd2532: data = 1'd0;
		12'd2533: data = 1'd0;
		12'd2534: data = 1'd0;
		12'd2535: data = 1'd1;
		12'd2536: data = 1'd1;
		12'd2537: data = 1'd1;
		12'd2538: data = 1'd1;
		12'd2539: data = 1'd0;
		12'd2540: data = 1'd0;
		12'd2541: data = 1'd1;
		12'd2542: data = 1'd0;
		12'd2543: data = 1'd0;
		12'd2544: data = 1'd0;
		12'd2545: data = 1'd0;
		12'd2546: data = 1'd0;
		12'd2547: data = 1'd0;
		12'd2548: data = 1'd0;
		12'd2549: data = 1'd0;
		12'd2550: data = 1'd0;
		12'd2551: data = 1'd0;
		12'd2552: data = 1'd1;
		12'd2553: data = 1'd1;
		12'd2554: data = 1'd1;
		12'd2555: data = 1'd1;
		12'd2556: data = 1'd1;
		12'd2557: data = 1'd1;
		12'd2558: data = 1'd0;
		12'd2559: data = 1'd0;
		12'd2560: data = 1'd0;
		12'd2561: data = 1'd0;
		12'd2562: data = 1'd0;
		12'd2563: data = 1'd0;
		12'd2564: data = 1'd0;
		12'd2565: data = 1'd0;
		12'd2566: data = 1'd0;
		12'd2567: data = 1'd0;
		12'd2568: data = 1'd0;
		12'd2569: data = 1'd0;
		12'd2570: data = 1'd0;
		12'd2571: data = 1'd0;
		12'd2572: data = 1'd0;
		12'd2573: data = 1'd0;
		12'd2574: data = 1'd1;
		12'd2575: data = 1'd0;
		12'd2576: data = 1'd1;
		12'd2577: data = 1'd0;
		12'd2578: data = 1'd0;
		12'd2579: data = 1'd0;
		12'd2580: data = 1'd0;
		12'd2581: data = 1'd0;
		12'd2582: data = 1'd0;
		12'd2583: data = 1'd0;
		12'd2584: data = 1'd0;
		12'd2585: data = 1'd0;
		12'd2586: data = 1'd0;
		12'd2587: data = 1'd0;
		12'd2588: data = 1'd0;
		12'd2589: data = 1'd1;
		12'd2590: data = 1'd0;
		12'd2591: data = 1'd1;
		12'd2592: data = 1'd0;
		12'd2593: data = 1'd1;
		12'd2594: data = 1'd0;
		12'd2595: data = 1'd0;
		12'd2596: data = 1'd0;
		12'd2597: data = 1'd0;
		12'd2598: data = 1'd0;
		12'd2599: data = 1'd0;
		12'd2600: data = 1'd0;
		12'd2601: data = 1'd0;
		12'd2602: data = 1'd0;
		12'd2603: data = 1'd0;
		12'd2604: data = 1'd1;
		12'd2605: data = 1'd0;
		12'd2606: data = 1'd1;
		12'd2607: data = 1'd0;
		12'd2608: data = 1'd0;
		12'd2609: data = 1'd1;
		12'd2610: data = 1'd0;
		12'd2611: data = 1'd0;
		12'd2612: data = 1'd0;
		12'd2613: data = 1'd0;
		12'd2614: data = 1'd0;
		12'd2615: data = 1'd0;
		12'd2616: data = 1'd0;
		12'd2617: data = 1'd0;
		12'd2618: data = 1'd0;
		12'd2619: data = 1'd1;
		12'd2620: data = 1'd0;
		12'd2621: data = 1'd1;
		12'd2622: data = 1'd0;
		12'd2623: data = 1'd1;
		12'd2624: data = 1'd0;
		12'd2625: data = 1'd0;
		12'd2626: data = 1'd1;
		12'd2627: data = 1'd1;
		12'd2628: data = 1'd0;
		12'd2629: data = 1'd0;
		12'd2630: data = 1'd1;
		12'd2631: data = 1'd1;
		12'd2632: data = 1'd0;
		12'd2633: data = 1'd1;
		12'd2634: data = 1'd1;
		12'd2635: data = 1'd0;
		12'd2636: data = 1'd0;
		12'd2637: data = 1'd1;
		12'd2638: data = 1'd0;
		12'd2639: data = 1'd1;
		12'd2640: data = 1'd0;
		12'd2641: data = 1'd0;
		12'd2642: data = 1'd1;
		12'd2643: data = 1'd0;
		12'd2644: data = 1'd0;
		12'd2645: data = 1'd1;
		12'd2646: data = 1'd0;
		12'd2647: data = 1'd1;
		12'd2648: data = 1'd0;
		12'd2649: data = 1'd0;
		12'd2650: data = 1'd0;
		12'd2651: data = 1'd0;
		12'd2652: data = 1'd1;
		12'd2653: data = 1'd0;
		12'd2654: data = 1'd1;
		12'd2655: data = 1'd0;
		12'd2656: data = 1'd0;
		12'd2657: data = 1'd0;
		12'd2658: data = 1'd1;
		12'd2659: data = 1'd0;
		12'd2660: data = 1'd1;
		12'd2661: data = 1'd1;
		12'd2662: data = 1'd0;
		12'd2663: data = 1'd1;
		12'd2664: data = 1'd1;
		12'd2665: data = 1'd0;
		12'd2666: data = 1'd1;
		12'd2667: data = 1'd0;
		12'd2668: data = 1'd0;
		12'd2669: data = 1'd1;
		12'd2670: data = 1'd0;
		12'd2671: data = 1'd0;
		12'd2672: data = 1'd0;
		12'd2673: data = 1'd0;
		12'd2674: data = 1'd0;
		12'd2675: data = 1'd1;
		12'd2676: data = 1'd1;
		12'd2677: data = 1'd1;
		12'd2678: data = 1'd1;
		12'd2679: data = 1'd0;
		12'd2680: data = 1'd1;
		12'd2681: data = 1'd0;
		12'd2682: data = 1'd1;
		12'd2683: data = 1'd1;
		12'd2684: data = 1'd1;
		12'd2685: data = 1'd0;
		12'd2686: data = 1'd0;
		12'd2687: data = 1'd1;
		12'd2688: data = 1'd0;
		12'd2689: data = 1'd0;
		12'd2690: data = 1'd0;
		12'd2691: data = 1'd1;
		12'd2692: data = 1'd1;
		12'd2693: data = 1'd0;
		12'd2694: data = 1'd1;
		12'd2695: data = 1'd0;
		12'd2696: data = 1'd1;
		12'd2697: data = 1'd0;
		12'd2698: data = 1'd0;
		12'd2699: data = 1'd1;
		12'd2700: data = 1'd0;
		12'd2701: data = 1'd1;
		12'd2702: data = 1'd1;
		12'd2703: data = 1'd0;
		12'd2704: data = 1'd0;
		12'd2705: data = 1'd0;
		12'd2706: data = 1'd0;
		12'd2707: data = 1'd0;
		12'd2708: data = 1'd0;
		12'd2709: data = 1'd0;
		12'd2710: data = 1'd1;
		12'd2711: data = 1'd1;
		12'd2712: data = 1'd0;
		12'd2713: data = 1'd1;
		12'd2714: data = 1'd0;
		12'd2715: data = 1'd1;
		12'd2716: data = 1'd0;
		12'd2717: data = 1'd0;
		12'd2718: data = 1'd0;
		12'd2719: data = 1'd1;
		12'd2720: data = 1'd0;
		12'd2721: data = 1'd0;
		12'd2722: data = 1'd0;
		12'd2723: data = 1'd0;
		12'd2724: data = 1'd0;
		12'd2725: data = 1'd0;
		12'd2726: data = 1'd0;
		12'd2727: data = 1'd1;
		12'd2728: data = 1'd0;
		12'd2729: data = 1'd1;
		12'd2730: data = 1'd0;
		12'd2731: data = 1'd1;
		12'd2732: data = 1'd1;
		12'd2733: data = 1'd0;
		12'd2734: data = 1'd1;
		12'd2735: data = 1'd0;
		12'd2736: data = 1'd0;
		12'd2737: data = 1'd0;
		12'd2738: data = 1'd0;
		12'd2739: data = 1'd0;
		12'd2740: data = 1'd1;
		12'd2741: data = 1'd1;
		12'd2742: data = 1'd1;
		12'd2743: data = 1'd1;
		12'd2744: data = 1'd0;
		12'd2745: data = 1'd1;
		12'd2746: data = 1'd1;
		12'd2747: data = 1'd0;
		12'd2748: data = 1'd1;
		12'd2749: data = 1'd0;
		12'd2750: data = 1'd1;
		12'd2751: data = 1'd1;
		12'd2752: data = 1'd0;
		12'd2753: data = 1'd0;
		12'd2754: data = 1'd0;
		12'd2755: data = 1'd0;
		12'd2756: data = 1'd1;
		12'd2757: data = 1'd1;
		12'd2758: data = 1'd1;
		12'd2759: data = 1'd1;
		12'd2760: data = 1'd0;
		12'd2761: data = 1'd1;
		12'd2762: data = 1'd0;
		12'd2763: data = 1'd0;
		12'd2764: data = 1'd1;
		12'd2765: data = 1'd0;
		12'd2766: data = 1'd1;
		12'd2767: data = 1'd0;
		12'd2768: data = 1'd0;
		12'd2769: data = 1'd0;
		12'd2770: data = 1'd0;
		12'd2771: data = 1'd0;
		12'd2772: data = 1'd0;
		12'd2773: data = 1'd0;
		12'd2774: data = 1'd0;
		12'd2775: data = 1'd0;
		12'd2776: data = 1'd1;
		12'd2777: data = 1'd1;
		12'd2778: data = 1'd0;
		12'd2779: data = 1'd1;
		12'd2780: data = 1'd0;
		12'd2781: data = 1'd1;
		12'd2782: data = 1'd0;
		12'd2783: data = 1'd0;
		12'd2784: data = 1'd0;
		12'd2785: data = 1'd0;
		12'd2786: data = 1'd0;
		12'd2787: data = 1'd0;
		12'd2788: data = 1'd0;
		12'd2789: data = 1'd1;
		12'd2790: data = 1'd0;
		12'd2791: data = 1'd0;
		12'd2792: data = 1'd0;
		12'd2793: data = 1'd1;
		12'd2794: data = 1'd1;
		12'd2795: data = 1'd0;
		12'd2796: data = 1'd0;
		12'd2797: data = 1'd1;
		12'd2798: data = 1'd0;
		12'd2799: data = 1'd1;
		12'd2800: data = 1'd0;
		12'd2801: data = 1'd0;
		12'd2802: data = 1'd0;
		12'd2803: data = 1'd0;
		12'd2804: data = 1'd0;
		12'd2805: data = 1'd0;
		12'd2806: data = 1'd1;
		12'd2807: data = 1'd1;
		12'd2808: data = 1'd0;
		12'd2809: data = 1'd0;
		12'd2810: data = 1'd0;
		12'd2811: data = 1'd0;
		12'd2812: data = 1'd1;
		12'd2813: data = 1'd0;
		12'd2814: data = 1'd1;
		12'd2815: data = 1'd0;
		12'd2816: data = 1'd0;
		12'd2817: data = 1'd1;
		12'd2818: data = 1'd0;
		12'd2819: data = 1'd0;
		12'd2820: data = 1'd0;
		12'd2821: data = 1'd0;
		12'd2822: data = 1'd0;
		12'd2823: data = 1'd0;
		12'd2824: data = 1'd0;
		12'd2825: data = 1'd0;
		12'd2826: data = 1'd0;
		12'd2827: data = 1'd0;
		12'd2828: data = 1'd0;
		12'd2829: data = 1'd1;
		12'd2830: data = 1'd0;
		12'd2831: data = 1'd0;
		12'd2832: data = 1'd0;
		12'd2833: data = 1'd1;
		12'd2834: data = 1'd0;
		12'd2835: data = 1'd0;
		12'd2836: data = 1'd0;
		12'd2837: data = 1'd0;
		12'd2838: data = 1'd0;
		12'd2839: data = 1'd0;
		12'd2840: data = 1'd0;
		12'd2841: data = 1'd0;
		12'd2842: data = 1'd0;
		12'd2843: data = 1'd0;
		12'd2844: data = 1'd1;
		12'd2845: data = 1'd0;
		12'd2846: data = 1'd0;
		12'd2847: data = 1'd1;
		12'd2848: data = 1'd1;
		12'd2849: data = 1'd0;
		12'd2850: data = 1'd1;
		12'd2851: data = 1'd0;
		12'd2852: data = 1'd0;
		12'd2853: data = 1'd0;
		12'd2854: data = 1'd0;
		12'd2855: data = 1'd0;
		12'd2856: data = 1'd0;
		12'd2857: data = 1'd0;
		12'd2858: data = 1'd0;
		12'd2859: data = 1'd1;
		12'd2860: data = 1'd0;
		12'd2861: data = 1'd0;
		12'd2862: data = 1'd1;
		12'd2863: data = 1'd0;
		12'd2864: data = 1'd1;
		12'd2865: data = 1'd0;
		12'd2866: data = 1'd1;
		12'd2867: data = 1'd0;
		12'd2868: data = 1'd1;
		12'd2869: data = 1'd0;
		12'd2870: data = 1'd1;
		12'd2871: data = 1'd0;
		12'd2872: data = 1'd1;
		12'd2873: data = 1'd0;
		12'd2874: data = 1'd0;
		12'd2875: data = 1'd0;
		12'd2876: data = 1'd0;
		12'd2877: data = 1'd1;
		12'd2878: data = 1'd0;
		12'd2879: data = 1'd1;
		12'd2880: data = 1'd1;
		12'd2881: data = 1'd1;
		12'd2882: data = 1'd1;
		12'd2883: data = 1'd0;
		12'd2884: data = 1'd1;
		12'd2885: data = 1'd0;
		12'd2886: data = 1'd0;
		12'd2887: data = 1'd1;
		12'd2888: data = 1'd0;
		12'd2889: data = 1'd0;
		12'd2890: data = 1'd0;
		12'd2891: data = 1'd1;
		12'd2892: data = 1'd0;
		12'd2893: data = 1'd1;
		12'd2894: data = 1'd0;
		12'd2895: data = 1'd1;
		12'd2896: data = 1'd1;
		12'd2897: data = 1'd1;
		12'd2898: data = 1'd0;
		12'd2899: data = 1'd1;
		12'd2900: data = 1'd0;
		12'd2901: data = 1'd1;
		12'd2902: data = 1'd0;
		12'd2903: data = 1'd1;
		12'd2904: data = 1'd0;
		12'd2905: data = 1'd1;
		12'd2906: data = 1'd0;
		12'd2907: data = 1'd0;
		12'd2908: data = 1'd1;
		12'd2909: data = 1'd1;
		12'd2910: data = 1'd1;
		12'd2911: data = 1'd0;
		12'd2912: data = 1'd1;
		12'd2913: data = 1'd1;
		12'd2914: data = 1'd0;
		12'd2915: data = 1'd1;
		12'd2916: data = 1'd0;
		12'd2917: data = 1'd1;
		12'd2918: data = 1'd0;
		12'd2919: data = 1'd0;
		12'd2920: data = 1'd1;
		12'd2921: data = 1'd0;
		12'd2922: data = 1'd1;
		12'd2923: data = 1'd0;
		12'd2924: data = 1'd1;
		12'd2925: data = 1'd0;
		12'd2926: data = 1'd0;
		12'd2927: data = 1'd0;
		12'd2928: data = 1'd0;
		12'd2929: data = 1'd1;
		12'd2930: data = 1'd1;
		12'd2931: data = 1'd0;
		12'd2932: data = 1'd1;
		12'd2933: data = 1'd0;
		12'd2934: data = 1'd1;
		12'd2935: data = 1'd0;
		12'd2936: data = 1'd1;
		12'd2937: data = 1'd0;
		12'd2938: data = 1'd1;
		12'd2939: data = 1'd0;
		12'd2940: data = 1'd1;
		12'd2941: data = 1'd0;
		12'd2942: data = 1'd1;
		12'd2943: data = 1'd1;
		12'd2944: data = 1'd0;
		12'd2945: data = 1'd1;
		12'd2946: data = 1'd1;
		12'd2947: data = 1'd0;
		12'd2948: data = 1'd1;
		12'd2949: data = 1'd0;
		12'd2950: data = 1'd1;
		12'd2951: data = 1'd0;
		12'd2952: data = 1'd1;
		12'd2953: data = 1'd1;
		12'd2954: data = 1'd0;
		12'd2955: data = 1'd1;
		12'd2956: data = 1'd0;
		12'd2957: data = 1'd1;
		12'd2958: data = 1'd0;
		12'd2959: data = 1'd1;
		12'd2960: data = 1'd1;
		12'd2961: data = 1'd0;
		12'd2962: data = 1'd1;
		12'd2963: data = 1'd0;
		12'd2964: data = 1'd1;
		12'd2965: data = 1'd1;
		12'd2966: data = 1'd0;
		12'd2967: data = 1'd1;
		12'd2968: data = 1'd0;
		12'd2969: data = 1'd1;
		12'd2970: data = 1'd0;
		12'd2971: data = 1'd1;
		12'd2972: data = 1'd0;
		12'd2973: data = 1'd1;
		12'd2974: data = 1'd0;
		12'd2975: data = 1'd1;
		12'd2976: data = 1'd1;
		12'd2977: data = 1'd0;
		12'd2978: data = 1'd1;
		12'd2979: data = 1'd1;
		12'd2980: data = 1'd0;
		12'd2981: data = 1'd1;
		12'd2982: data = 1'd0;
		12'd2983: data = 1'd1;
		12'd2984: data = 1'd0;
		12'd2985: data = 1'd1;
		12'd2986: data = 1'd1;
		12'd2987: data = 1'd0;
		12'd2988: data = 1'd1;
		12'd2989: data = 1'd0;
		12'd2990: data = 1'd1;
		12'd2991: data = 1'd0;
		12'd2992: data = 1'd1;
		12'd2993: data = 1'd0;
		12'd2994: data = 1'd0;
		12'd2995: data = 1'd0;
		12'd2996: data = 1'd0;
		12'd2997: data = 1'd1;
		12'd2998: data = 1'd0;
		12'd2999: data = 1'd0;
		12'd3000: data = 1'd1;
		12'd3001: data = 1'd0;
		12'd3002: data = 1'd1;
		12'd3003: data = 1'd0;
		12'd3004: data = 1'd1;
		12'd3005: data = 1'd0;
		12'd3006: data = 1'd1;
		12'd3007: data = 1'd0;
		12'd3008: data = 1'd1;
		12'd3009: data = 1'd1;
		12'd3010: data = 1'd0;
		12'd3011: data = 1'd0;
		12'd3012: data = 1'd1;
		12'd3013: data = 1'd1;
		12'd3014: data = 1'd0;
		12'd3015: data = 1'd1;
		12'd3016: data = 1'd1;
		12'd3017: data = 1'd0;
		12'd3018: data = 1'd1;
		12'd3019: data = 1'd0;
		12'd3020: data = 1'd0;
		12'd3021: data = 1'd1;
		12'd3022: data = 1'd0;
		12'd3023: data = 1'd1;
		12'd3024: data = 1'd0;
		12'd3025: data = 1'd1;
		12'd3026: data = 1'd0;
		12'd3027: data = 1'd0;
		12'd3028: data = 1'd1;
		12'd3029: data = 1'd0;
		12'd3030: data = 1'd0;
		12'd3031: data = 1'd1;
		12'd3032: data = 1'd0;
		12'd3033: data = 1'd1;
		12'd3034: data = 1'd1;
		12'd3035: data = 1'd0;
		12'd3036: data = 1'd1;
		12'd3037: data = 1'd0;
		12'd3038: data = 1'd0;
		12'd3039: data = 1'd1;
		12'd3040: data = 1'd0;
		12'd3041: data = 1'd0;
		12'd3042: data = 1'd1;
		12'd3043: data = 1'd1;
		12'd3044: data = 1'd1;
		12'd3045: data = 1'd0;
		12'd3046: data = 1'd1;
		12'd3047: data = 1'd1;
		12'd3048: data = 1'd0;
		12'd3049: data = 1'd1;
		12'd3050: data = 1'd0;
		12'd3051: data = 1'd0;
		12'd3052: data = 1'd1;
		12'd3053: data = 1'd0;
		12'd3054: data = 1'd1;
		12'd3055: data = 1'd0;
		12'd3056: data = 1'd0;
		12'd3057: data = 1'd0;
		12'd3058: data = 1'd0;
		12'd3059: data = 1'd0;
		12'd3060: data = 1'd1;
		12'd3061: data = 1'd1;
		12'd3062: data = 1'd1;
		12'd3063: data = 1'd0;
		12'd3064: data = 1'd1;
		12'd3065: data = 1'd1;
		12'd3066: data = 1'd0;
		12'd3067: data = 1'd1;
		12'd3068: data = 1'd0;
		12'd3069: data = 1'd1;
		12'd3070: data = 1'd0;
		12'd3071: data = 1'd1;
		12'd3072: data = 1'd0;
		12'd3073: data = 1'd1;
		12'd3074: data = 1'd0;
		12'd3075: data = 1'd0;
		12'd3076: data = 1'd0;
		12'd3077: data = 1'd0;
		12'd3078: data = 1'd0;
		12'd3079: data = 1'd0;
		12'd3080: data = 1'd0;
		12'd3081: data = 1'd0;
		12'd3082: data = 1'd0;
		12'd3083: data = 1'd0;
		12'd3084: data = 1'd1;
		12'd3085: data = 1'd0;
		12'd3086: data = 1'd0;
		12'd3087: data = 1'd1;
		12'd3088: data = 1'd1;
		12'd3089: data = 1'd0;
		12'd3090: data = 1'd1;
		12'd3091: data = 1'd0;
		12'd3092: data = 1'd1;
		12'd3093: data = 1'd0;
		12'd3094: data = 1'd1;
		12'd3095: data = 1'd1;
		12'd3096: data = 1'd0;
		12'd3097: data = 1'd0;
		12'd3098: data = 1'd0;
		12'd3099: data = 1'd0;
		12'd3100: data = 1'd1;
		12'd3101: data = 1'd0;
		12'd3102: data = 1'd1;
		12'd3103: data = 1'd1;
		12'd3104: data = 1'd1;
		12'd3105: data = 1'd0;
		12'd3106: data = 1'd1;
		12'd3107: data = 1'd0;
		12'd3108: data = 1'd1;
		12'd3109: data = 1'd0;
		12'd3110: data = 1'd1;
		12'd3111: data = 1'd1;
		12'd3112: data = 1'd0;
		12'd3113: data = 1'd0;
		12'd3114: data = 1'd1;
		12'd3115: data = 1'd0;
		12'd3116: data = 1'd1;
		12'd3117: data = 1'd0;
		12'd3118: data = 1'd0;
		12'd3119: data = 1'd1;
		12'd3120: data = 1'd1;
		12'd3121: data = 1'd0;
		12'd3122: data = 1'd1;
		12'd3123: data = 1'd0;
		12'd3124: data = 1'd1;
		12'd3125: data = 1'd0;
		12'd3126: data = 1'd1;
		12'd3127: data = 1'd0;
		12'd3128: data = 1'd0;
		12'd3129: data = 1'd1;
		12'd3130: data = 1'd0;
		12'd3131: data = 1'd0;
		12'd3132: data = 1'd1;
		12'd3133: data = 1'd1;
		12'd3134: data = 1'd0;
		12'd3135: data = 1'd1;
		12'd3136: data = 1'd1;
		12'd3137: data = 1'd1;
		12'd3138: data = 1'd0;
		12'd3139: data = 1'd1;
		12'd3140: data = 1'd0;
		12'd3141: data = 1'd1;
		12'd3142: data = 1'd0;
		12'd3143: data = 1'd1;
		12'd3144: data = 1'd0;
		12'd3145: data = 1'd1;
		12'd3146: data = 1'd0;
		12'd3147: data = 1'd1;
		12'd3148: data = 1'd0;
		12'd3149: data = 1'd1;
		12'd3150: data = 1'd0;
		12'd3151: data = 1'd0;
		12'd3152: data = 1'd1;
		12'd3153: data = 1'd1;
		12'd3154: data = 1'd0;
		12'd3155: data = 1'd1;
		12'd3156: data = 1'd0;
		12'd3157: data = 1'd1;
		12'd3158: data = 1'd0;
		12'd3159: data = 1'd1;
		12'd3160: data = 1'd0;
		12'd3161: data = 1'd0;
		12'd3162: data = 1'd1;
		12'd3163: data = 1'd0;
		12'd3164: data = 1'd1;
		12'd3165: data = 1'd0;
		12'd3166: data = 1'd1;
		12'd3167: data = 1'd0;
		12'd3168: data = 1'd0;
		12'd3169: data = 1'd1;
		12'd3170: data = 1'd1;
		12'd3171: data = 1'd1;
		12'd3172: data = 1'd0;
		12'd3173: data = 1'd0;
		12'd3174: data = 1'd1;
		12'd3175: data = 1'd0;
		12'd3176: data = 1'd1;
		12'd3177: data = 1'd0;
		12'd3178: data = 1'd1;
		12'd3179: data = 1'd0;
		12'd3180: data = 1'd1;
		12'd3181: data = 1'd0;
		12'd3182: data = 1'd1;
		12'd3183: data = 1'd0;
		12'd3184: data = 1'd0;
		12'd3185: data = 1'd1;
		12'd3186: data = 1'd1;
		12'd3187: data = 1'd0;
		12'd3188: data = 1'd1;
		12'd3189: data = 1'd0;
		12'd3190: data = 1'd1;
		12'd3191: data = 1'd0;
		12'd3192: data = 1'd1;
		12'd3193: data = 1'd0;
		12'd3194: data = 1'd0;
		12'd3195: data = 1'd1;
		12'd3196: data = 1'd0;
		12'd3197: data = 1'd1;
		12'd3198: data = 1'd0;
		12'd3199: data = 1'd1;
		12'd3200: data = 1'd0;
		12'd3201: data = 1'd0;
		12'd3202: data = 1'd1;
		12'd3203: data = 1'd0;
		12'd3204: data = 1'd1;
		12'd3205: data = 1'd0;
		12'd3206: data = 1'd0;
		12'd3207: data = 1'd1;
		12'd3208: data = 1'd0;
		12'd3209: data = 1'd1;
		12'd3210: data = 1'd0;
		12'd3211: data = 1'd1;
		12'd3212: data = 1'd0;
		12'd3213: data = 1'd1;
		12'd3214: data = 1'd0;
		12'd3215: data = 1'd1;
		12'd3216: data = 1'd1;
		12'd3217: data = 1'd0;
		12'd3218: data = 1'd1;
		12'd3219: data = 1'd1;
		12'd3220: data = 1'd0;
		12'd3221: data = 1'd1;
		12'd3222: data = 1'd0;
		12'd3223: data = 1'd1;
		12'd3224: data = 1'd0;
		12'd3225: data = 1'd1;
		12'd3226: data = 1'd0;
		12'd3227: data = 1'd1;
		12'd3228: data = 1'd1;
		12'd3229: data = 1'd0;
		12'd3230: data = 1'd1;
		12'd3231: data = 1'd0;
		12'd3232: data = 1'd1;
		12'd3233: data = 1'd1;
		12'd3234: data = 1'd0;
		12'd3235: data = 1'd1;
		12'd3236: data = 1'd0;
		12'd3237: data = 1'd1;
		12'd3238: data = 1'd0;
		12'd3239: data = 1'd1;
		12'd3240: data = 1'd1;
		12'd3241: data = 1'd0;
		12'd3242: data = 1'd1;
		12'd3243: data = 1'd0;
		12'd3244: data = 1'd1;
		12'd3245: data = 1'd0;
		12'd3246: data = 1'd1;
		12'd3247: data = 1'd0;
		12'd3248: data = 1'd1;
		12'd3249: data = 1'd1;
		12'd3250: data = 1'd0;
		12'd3251: data = 1'd1;
		12'd3252: data = 1'd1;
		12'd3253: data = 1'd0;
		12'd3254: data = 1'd1;
		12'd3255: data = 1'd0;
		12'd3256: data = 1'd1;
		12'd3257: data = 1'd0;
		12'd3258: data = 1'd1;
		12'd3259: data = 1'd0;
		12'd3260: data = 1'd1;
		12'd3261: data = 1'd1;
		12'd3262: data = 1'd0;
		12'd3263: data = 1'd1;
		12'd3264: data = 1'd1;
		12'd3265: data = 1'd1;
		12'd3266: data = 1'd0;
		12'd3267: data = 1'd0;
		12'd3268: data = 1'd0;
		12'd3269: data = 1'd0;
		12'd3270: data = 1'd1;
		12'd3271: data = 1'd0;
		12'd3272: data = 1'd1;
		12'd3273: data = 1'd1;
		12'd3274: data = 1'd0;
		12'd3275: data = 1'd1;
		12'd3276: data = 1'd0;
		12'd3277: data = 1'd1;
		12'd3278: data = 1'd0;
		12'd3279: data = 1'd1;
		12'd3280: data = 1'd1;
		12'd3281: data = 1'd1;
		12'd3282: data = 1'd1;
		12'd3283: data = 1'd0;
		12'd3284: data = 1'd0;
		12'd3285: data = 1'd1;
		12'd3286: data = 1'd1;
		12'd3287: data = 1'd0;
		12'd3288: data = 1'd1;
		12'd3289: data = 1'd0;
		12'd3290: data = 1'd0;
		12'd3291: data = 1'd1;
		12'd3292: data = 1'd0;
		12'd3293: data = 1'd1;
		12'd3294: data = 1'd0;
		12'd3295: data = 1'd1;
		12'd3296: data = 1'd1;
		12'd3297: data = 1'd1;
		12'd3298: data = 1'd1;
		12'd3299: data = 1'd0;
		12'd3300: data = 1'd0;
		12'd3301: data = 1'd1;
		12'd3302: data = 1'd0;
		12'd3303: data = 1'd1;
		12'd3304: data = 1'd1;
		12'd3305: data = 1'd0;
		12'd3306: data = 1'd1;
		12'd3307: data = 1'd0;
		12'd3308: data = 1'd0;
		12'd3309: data = 1'd1;
		12'd3310: data = 1'd0;
		12'd3311: data = 1'd1;
		12'd3312: data = 1'd1;
		12'd3313: data = 1'd1;
		12'd3314: data = 1'd1;
		12'd3315: data = 1'd0;
		12'd3316: data = 1'd0;
		12'd3317: data = 1'd1;
		12'd3318: data = 1'd0;
		12'd3319: data = 1'd1;
		12'd3320: data = 1'd0;
		12'd3321: data = 1'd1;
		12'd3322: data = 1'd1;
		12'd3323: data = 1'd0;
		12'd3324: data = 1'd1;
		12'd3325: data = 1'd0;
		12'd3326: data = 1'd1;
		12'd3327: data = 1'd0;
		12'd3328: data = 1'd1;
		12'd3329: data = 1'd0;
		12'd3330: data = 1'd1;
		12'd3331: data = 1'd1;
		12'd3332: data = 1'd0;
		12'd3333: data = 1'd0;
		12'd3334: data = 1'd1;
		12'd3335: data = 1'd0;
		12'd3336: data = 1'd0;
		12'd3337: data = 1'd1;
		12'd3338: data = 1'd0;
		12'd3339: data = 1'd1;
		12'd3340: data = 1'd0;
		12'd3341: data = 1'd1;
		12'd3342: data = 1'd0;
		12'd3343: data = 1'd0;
		12'd3344: data = 1'd1;
		12'd3345: data = 1'd0;
		12'd3346: data = 1'd1;
		12'd3347: data = 1'd0;
		12'd3348: data = 1'd1;
		12'd3349: data = 1'd0;
		12'd3350: data = 1'd1;
		12'd3351: data = 1'd0;
		12'd3352: data = 1'd1;
		12'd3353: data = 1'd0;
		12'd3354: data = 1'd0;
		12'd3355: data = 1'd1;
		12'd3356: data = 1'd1;
		12'd3357: data = 1'd0;
		12'd3358: data = 1'd1;
		12'd3359: data = 1'd0;
		12'd3360: data = 1'd0;
		12'd3361: data = 1'd0;
		12'd3362: data = 1'd1;
		12'd3363: data = 1'd0;
		12'd3364: data = 1'd1;
		12'd3365: data = 1'd0;
		12'd3366: data = 1'd1;
		12'd3367: data = 1'd0;
		12'd3368: data = 1'd1;
		12'd3369: data = 1'd1;
		12'd3370: data = 1'd0;
		12'd3371: data = 1'd1;
		12'd3372: data = 1'd0;
		12'd3373: data = 1'd0;
		12'd3374: data = 1'd1;
		12'd3375: data = 1'd0;
		12'd3376: data = 1'd1;
		12'd3377: data = 1'd1;
		12'd3378: data = 1'd0;
		12'd3379: data = 1'd1;
		12'd3380: data = 1'd0;
		12'd3381: data = 1'd1;
		12'd3382: data = 1'd0;
		12'd3383: data = 1'd1;
		12'd3384: data = 1'd0;
		12'd3385: data = 1'd1;
		12'd3386: data = 1'd0;
		12'd3387: data = 1'd1;
		12'd3388: data = 1'd0;
		12'd3389: data = 1'd1;
		12'd3390: data = 1'd0;
		12'd3391: data = 1'd1;
		12'd3392: data = 1'd1;
		12'd3393: data = 1'd1;
		12'd3394: data = 1'd0;
		12'd3395: data = 1'd1;
		12'd3396: data = 1'd0;
		12'd3397: data = 1'd1;
		12'd3398: data = 1'd0;
		12'd3399: data = 1'd1;
		12'd3400: data = 1'd0;
		12'd3401: data = 1'd1;
		12'd3402: data = 1'd0;
		12'd3403: data = 1'd0;
		12'd3404: data = 1'd1;
		12'd3405: data = 1'd0;
		12'd3406: data = 1'd1;
		12'd3407: data = 1'd0;
		12'd3408: data = 1'd0;
		12'd3409: data = 1'd1;
		12'd3410: data = 1'd1;
		12'd3411: data = 1'd1;
		12'd3412: data = 1'd0;
		12'd3413: data = 1'd1;
		12'd3414: data = 1'd0;
		12'd3415: data = 1'd0;
		12'd3416: data = 1'd1;
		12'd3417: data = 1'd0;
		12'd3418: data = 1'd1;
		12'd3419: data = 1'd0;
		12'd3420: data = 1'd1;
		12'd3421: data = 1'd0;
		12'd3422: data = 1'd1;
		12'd3423: data = 1'd0;
		12'd3424: data = 1'd0;
		12'd3425: data = 1'd1;
		12'd3426: data = 1'd1;
		12'd3427: data = 1'd0;
		12'd3428: data = 1'd1;
		12'd3429: data = 1'd0;
		12'd3430: data = 1'd1;
		12'd3431: data = 1'd0;
		12'd3432: data = 1'd1;
		12'd3433: data = 1'd0;
		12'd3434: data = 1'd1;
		12'd3435: data = 1'd0;
		12'd3436: data = 1'd0;
		12'd3437: data = 1'd1;
		12'd3438: data = 1'd0;
		12'd3439: data = 1'd1;
		12'd3440: data = 1'd0;
		12'd3441: data = 1'd0;
		12'd3442: data = 1'd1;
		12'd3443: data = 1'd0;
		12'd3444: data = 1'd1;
		12'd3445: data = 1'd0;
		12'd3446: data = 1'd1;
		12'd3447: data = 1'd0;
		12'd3448: data = 1'd0;
		12'd3449: data = 1'd1;
		12'd3450: data = 1'd0;
		12'd3451: data = 1'd1;
		12'd3452: data = 1'd0;
		12'd3453: data = 1'd1;
		12'd3454: data = 1'd0;
		12'd3455: data = 1'd1;
		12'd3456: data = 1'd1;
		12'd3457: data = 1'd0;
		12'd3458: data = 1'd1;
		12'd3459: data = 1'd1;
		12'd3460: data = 1'd0;
		12'd3461: data = 1'd1;
		12'd3462: data = 1'd0;
		12'd3463: data = 1'd1;
		12'd3464: data = 1'd0;
		12'd3465: data = 1'd1;
		12'd3466: data = 1'd0;
		12'd3467: data = 1'd1;
		12'd3468: data = 1'd0;
		12'd3469: data = 1'd0;
		12'd3470: data = 1'd1;
		12'd3471: data = 1'd0;
		12'd3472: data = 1'd1;
		12'd3473: data = 1'd0;
		12'd3474: data = 1'd0;
		12'd3475: data = 1'd1;
		12'd3476: data = 1'd0;
		12'd3477: data = 1'd1;
		12'd3478: data = 1'd0;
		12'd3479: data = 1'd1;
		12'd3480: data = 1'd0;
		12'd3481: data = 1'd0;
		12'd3482: data = 1'd1;
		12'd3483: data = 1'd0;
		12'd3484: data = 1'd1;
		12'd3485: data = 1'd0;
		12'd3486: data = 1'd1;
		12'd3487: data = 1'd0;
		12'd3488: data = 1'd1;
		12'd3489: data = 1'd1;
		12'd3490: data = 1'd0;
		12'd3491: data = 1'd1;
		12'd3492: data = 1'd0;
		12'd3493: data = 1'd0;
		12'd3494: data = 1'd1;
		12'd3495: data = 1'd0;
		12'd3496: data = 1'd1;
		12'd3497: data = 1'd0;
		12'd3498: data = 1'd1;
		12'd3499: data = 1'd0;
		12'd3500: data = 1'd1;
		12'd3501: data = 1'd0;
		12'd3502: data = 1'd1;
		12'd3503: data = 1'd0;
		12'd3504: data = 1'd1;
		12'd3505: data = 1'd1;
		12'd3506: data = 1'd0;
		12'd3507: data = 1'd0;
		12'd3508: data = 1'd1;
		12'd3509: data = 1'd0;
		12'd3510: data = 1'd1;
		12'd3511: data = 1'd0;
		12'd3512: data = 1'd1;
		12'd3513: data = 1'd0;
		12'd3514: data = 1'd1;
		12'd3515: data = 1'd1;
		12'd3516: data = 1'd0;
		12'd3517: data = 1'd1;
		12'd3518: data = 1'd0;
		12'd3519: data = 1'd1;
		12'd3520: data = 1'd1;
		12'd3521: data = 1'd1;
		12'd3522: data = 1'd1;
		12'd3523: data = 1'd0;
		12'd3524: data = 1'd0;
		12'd3525: data = 1'd0;
		12'd3526: data = 1'd1;
		12'd3527: data = 1'd1;
		12'd3528: data = 1'd0;
		12'd3529: data = 1'd1;
		12'd3530: data = 1'd0;
		12'd3531: data = 1'd1;
		12'd3532: data = 1'd0;
		12'd3533: data = 1'd1;
		12'd3534: data = 1'd0;
		12'd3535: data = 1'd1;
		12'd3536: data = 1'd1;
		12'd3537: data = 1'd1;
		12'd3538: data = 1'd1;
		12'd3539: data = 1'd0;
		12'd3540: data = 1'd0;
		12'd3541: data = 1'd0;
		12'd3542: data = 1'd1;
		12'd3543: data = 1'd1;
		12'd3544: data = 1'd0;
		12'd3545: data = 1'd1;
		12'd3546: data = 1'd0;
		12'd3547: data = 1'd1;
		12'd3548: data = 1'd0;
		12'd3549: data = 1'd1;
		12'd3550: data = 1'd1;
		12'd3551: data = 1'd0;
		12'd3552: data = 1'd1;
		12'd3553: data = 1'd1;
		12'd3554: data = 1'd1;
		12'd3555: data = 1'd0;
		12'd3556: data = 1'd0;
		12'd3557: data = 1'd0;
		12'd3558: data = 1'd1;
		12'd3559: data = 1'd0;
		12'd3560: data = 1'd0;
		12'd3561: data = 1'd1;
		12'd3562: data = 1'd0;
		12'd3563: data = 1'd1;
		12'd3564: data = 1'd1;
		12'd3565: data = 1'd0;
		12'd3566: data = 1'd1;
		12'd3567: data = 1'd0;
		12'd3568: data = 1'd1;
		12'd3569: data = 1'd1;
		12'd3570: data = 1'd1;
		12'd3571: data = 1'd0;
		12'd3572: data = 1'd0;
		12'd3573: data = 1'd1;
		12'd3574: data = 1'd1;
		12'd3575: data = 1'd0;
		12'd3576: data = 1'd1;
		12'd3577: data = 1'd0;
		12'd3578: data = 1'd0;
		12'd3579: data = 1'd1;
		12'd3580: data = 1'd0;
		12'd3581: data = 1'd1;
		12'd3582: data = 1'd0;
		12'd3583: data = 1'd0;
		12'd3584: data = 1'd1;
		12'd3585: data = 1'd0;
		12'd3586: data = 1'd1;
		12'd3587: data = 1'd0;
		12'd3588: data = 1'd1;
		12'd3589: data = 1'd0;
		12'd3590: data = 1'd1;
		12'd3591: data = 1'd0;
		12'd3592: data = 1'd1;
		12'd3593: data = 1'd0;
		12'd3594: data = 1'd1;
		12'd3595: data = 1'd0;
		12'd3596: data = 1'd0;
		12'd3597: data = 1'd1;
		12'd3598: data = 1'd0;
		12'd3599: data = 1'd1;
		12'd3600: data = 1'd1;
		12'd3601: data = 1'd0;
		12'd3602: data = 1'd1;
		12'd3603: data = 1'd0;
		12'd3604: data = 1'd1;
		12'd3605: data = 1'd0;
		12'd3606: data = 1'd1;
		12'd3607: data = 1'd0;
		12'd3608: data = 1'd1;
		12'd3609: data = 1'd0;
		12'd3610: data = 1'd1;
		12'd3611: data = 1'd1;
		12'd3612: data = 1'd0;
		12'd3613: data = 1'd1;
		12'd3614: data = 1'd0;
		12'd3615: data = 1'd1;
		12'd3616: data = 1'd1;
		12'd3617: data = 1'd1;
		12'd3618: data = 1'd0;
		12'd3619: data = 1'd1;
		12'd3620: data = 1'd1;
		12'd3621: data = 1'd0;
		12'd3622: data = 1'd1;
		12'd3623: data = 1'd1;
		12'd3624: data = 1'd0;
		12'd3625: data = 1'd1;
		12'd3626: data = 1'd0;
		12'd3627: data = 1'd1;
		12'd3628: data = 1'd0;
		12'd3629: data = 1'd1;
		12'd3630: data = 1'd0;
		12'd3631: data = 1'd1;
		12'd3632: data = 1'd1;
		12'd3633: data = 1'd1;
		12'd3634: data = 1'd0;
		12'd3635: data = 1'd1;
		12'd3636: data = 1'd0;
		12'd3637: data = 1'd1;
		12'd3638: data = 1'd0;
		12'd3639: data = 1'd1;
		12'd3640: data = 1'd0;
		12'd3641: data = 1'd1;
		12'd3642: data = 1'd0;
		12'd3643: data = 1'd1;
		12'd3644: data = 1'd1;
		12'd3645: data = 1'd0;
		12'd3646: data = 1'd1;
		12'd3647: data = 1'd0;
		12'd3648: data = 1'd1;
		12'd3649: data = 1'd1;
		12'd3650: data = 1'd0;
		12'd3651: data = 1'd1;
		12'd3652: data = 1'd0;
		12'd3653: data = 1'd1;
		12'd3654: data = 1'd0;
		12'd3655: data = 1'd1;
		12'd3656: data = 1'd1;
		12'd3657: data = 1'd0;
		12'd3658: data = 1'd1;
		12'd3659: data = 1'd0;
		12'd3660: data = 1'd1;
		12'd3661: data = 1'd0;
		12'd3662: data = 1'd1;
		12'd3663: data = 1'd0;
		12'd3664: data = 1'd0;
		12'd3665: data = 1'd1;
		12'd3666: data = 1'd1;
		12'd3667: data = 1'd0;
		12'd3668: data = 1'd1;
		12'd3669: data = 1'd0;
		12'd3670: data = 1'd1;
		12'd3671: data = 1'd0;
		12'd3672: data = 1'd1;
		12'd3673: data = 1'd0;
		12'd3674: data = 1'd1;
		12'd3675: data = 1'd0;
		12'd3676: data = 1'd1;
		12'd3677: data = 1'd0;
		12'd3678: data = 1'd0;
		12'd3679: data = 1'd0;
		12'd3680: data = 1'd0;
		12'd3681: data = 1'd1;
		12'd3682: data = 1'd1;
		12'd3683: data = 1'd0;
		12'd3684: data = 1'd1;
		12'd3685: data = 1'd0;
		12'd3686: data = 1'd1;
		12'd3687: data = 1'd0;
		12'd3688: data = 1'd1;
		12'd3689: data = 1'd0;
		12'd3690: data = 1'd0;
		12'd3691: data = 1'd1;
		12'd3692: data = 1'd0;
		12'd3693: data = 1'd1;
		12'd3694: data = 1'd0;
		12'd3695: data = 1'd1;
		12'd3696: data = 1'd1;
		12'd3697: data = 1'd0;
		12'd3698: data = 1'd1;
		12'd3699: data = 1'd1;
		12'd3700: data = 1'd1;
		12'd3701: data = 1'd0;
		12'd3702: data = 1'd0;
		12'd3703: data = 1'd1;
		12'd3704: data = 1'd0;
		12'd3705: data = 1'd1;
		12'd3706: data = 1'd0;
		12'd3707: data = 1'd1;
		12'd3708: data = 1'd0;
		12'd3709: data = 1'd1;
		12'd3710: data = 1'd0;
		12'd3711: data = 1'd1;
		12'd3712: data = 1'd1;
		12'd3713: data = 1'd0;
		12'd3714: data = 1'd1;
		12'd3715: data = 1'd1;
		12'd3716: data = 1'd0;
		12'd3717: data = 1'd1;
		12'd3718: data = 1'd0;
		12'd3719: data = 1'd1;
		12'd3720: data = 1'd0;
		12'd3721: data = 1'd1;
		12'd3722: data = 1'd0;
		12'd3723: data = 1'd0;
		12'd3724: data = 1'd1;
		12'd3725: data = 1'd0;
		12'd3726: data = 1'd1;
		12'd3727: data = 1'd0;
		12'd3728: data = 1'd1;
		12'd3729: data = 1'd1;
		12'd3730: data = 1'd0;
		12'd3731: data = 1'd1;
		12'd3732: data = 1'd0;
		12'd3733: data = 1'd1;
		12'd3734: data = 1'd0;
		12'd3735: data = 1'd0;
		12'd3736: data = 1'd1;
		12'd3737: data = 1'd0;
		12'd3738: data = 1'd1;
		12'd3739: data = 1'd0;
		12'd3740: data = 1'd1;
		12'd3741: data = 1'd0;
		12'd3742: data = 1'd1;
		12'd3743: data = 1'd0;
		12'd3744: data = 1'd1;
		12'd3745: data = 1'd1;
		12'd3746: data = 1'd0;
		12'd3747: data = 1'd1;
		12'd3748: data = 1'd1;
		12'd3749: data = 1'd0;
		12'd3750: data = 1'd1;
		12'd3751: data = 1'd0;
		12'd3752: data = 1'd1;
		12'd3753: data = 1'd0;
		12'd3754: data = 1'd1;
		12'd3755: data = 1'd0;
		12'd3756: data = 1'd0;
		12'd3757: data = 1'd1;
		12'd3758: data = 1'd0;
		12'd3759: data = 1'd1;
		12'd3760: data = 1'd1;
		12'd3761: data = 1'd1;
		12'd3762: data = 1'd1;
		12'd3763: data = 1'd0;
		12'd3764: data = 1'd1;
		12'd3765: data = 1'd0;
		12'd3766: data = 1'd1;
		12'd3767: data = 1'd0;
		12'd3768: data = 1'd0;
		12'd3769: data = 1'd1;
		12'd3770: data = 1'd0;
		12'd3771: data = 1'd1;
		12'd3772: data = 1'd0;
		12'd3773: data = 1'd1;
		12'd3774: data = 1'd0;
		12'd3775: data = 1'd1;
		12'd3776: data = 1'd1;
		12'd3777: data = 1'd1;
		12'd3778: data = 1'd1;
		12'd3779: data = 1'd0;
		12'd3780: data = 1'd0;
		12'd3781: data = 1'd0;
		12'd3782: data = 1'd0;
		12'd3783: data = 1'd1;
		12'd3784: data = 1'd0;
		12'd3785: data = 1'd1;
		12'd3786: data = 1'd0;
		12'd3787: data = 1'd1;
		12'd3788: data = 1'd0;
		12'd3789: data = 1'd1;
		12'd3790: data = 1'd1;
		12'd3791: data = 1'd0;
		12'd3792: data = 1'd1;
		12'd3793: data = 1'd1;
		12'd3794: data = 1'd1;
		12'd3795: data = 1'd1;
		12'd3796: data = 1'd0;
		12'd3797: data = 1'd0;
		12'd3798: data = 1'd0;
		12'd3799: data = 1'd1;
		12'd3800: data = 1'd0;
		12'd3801: data = 1'd1;
		12'd3802: data = 1'd1;
		12'd3803: data = 1'd0;
		12'd3804: data = 1'd1;
		12'd3805: data = 1'd0;
		12'd3806: data = 1'd1;
		12'd3807: data = 1'd0;
		12'd3808: data = 1'd1;
		12'd3809: data = 1'd1;
		12'd3810: data = 1'd1;
		12'd3811: data = 1'd1;
		12'd3812: data = 1'd0;
		12'd3813: data = 1'd0;
		12'd3814: data = 1'd0;
		12'd3815: data = 1'd1;
		12'd3816: data = 1'd0;
		12'd3817: data = 1'd0;
		12'd3818: data = 1'd1;
		12'd3819: data = 1'd0;
		12'd3820: data = 1'd1;
		12'd3821: data = 1'd0;
		12'd3822: data = 1'd1;
		12'd3823: data = 1'd0;
		12'd3824: data = 1'd1;
		12'd3825: data = 1'd1;
		12'd3826: data = 1'd1;
		12'd3827: data = 1'd1;
		12'd3828: data = 1'd1;
		12'd3829: data = 1'd1;
		12'd3830: data = 1'd1;
		12'd3831: data = 1'd1;
		12'd3832: data = 1'd0;
		12'd3833: data = 1'd1;
		12'd3834: data = 1'd0;
		12'd3835: data = 1'd0;
		12'd3836: data = 1'd1;
		12'd3837: data = 1'd0;
		12'd3838: data = 1'd1;
		12'd3839: data = 1'd0;
		12'd3840: data = 1'd1;
		12'd3841: data = 1'd0;
		12'd3842: data = 1'd1;
		12'd3843: data = 1'd0;
		12'd3844: data = 1'd1;
		12'd3845: data = 1'd0;
		12'd3846: data = 1'd1;
		12'd3847: data = 1'd0;
		12'd3848: data = 1'd1;
		12'd3849: data = 1'd0;
		12'd3850: data = 1'd1;
		12'd3851: data = 1'd0;
		12'd3852: data = 1'd0;
		12'd3853: data = 1'd1;
		12'd3854: data = 1'd1;
		12'd3855: data = 1'd1;
		12'd3856: data = 1'd0;
		12'd3857: data = 1'd1;
		12'd3858: data = 1'd0;
		12'd3859: data = 1'd1;
		12'd3860: data = 1'd1;
		12'd3861: data = 1'd0;
		12'd3862: data = 1'd1;
		12'd3863: data = 1'd0;
		12'd3864: data = 1'd0;
		12'd3865: data = 1'd1;
		12'd3866: data = 1'd0;
		12'd3867: data = 1'd1;
		12'd3868: data = 1'd0;
		12'd3869: data = 1'd1;
		12'd3870: data = 1'd0;
		12'd3871: data = 1'd1;
		12'd3872: data = 1'd1;
		12'd3873: data = 1'd1;
		12'd3874: data = 1'd0;
		12'd3875: data = 1'd1;
		12'd3876: data = 1'd0;
		12'd3877: data = 1'd1;
		12'd3878: data = 1'd0;
		12'd3879: data = 1'd1;
		12'd3880: data = 1'd0;
		12'd3881: data = 1'd1;
		12'd3882: data = 1'd0;
		12'd3883: data = 1'd1;
		12'd3884: data = 1'd0;
		12'd3885: data = 1'd1;
		12'd3886: data = 1'd0;
		12'd3887: data = 1'd1;
		12'd3888: data = 1'd1;
		12'd3889: data = 1'd0;
		12'd3890: data = 1'd0;
		12'd3891: data = 1'd1;
		12'd3892: data = 1'd0;
		12'd3893: data = 1'd1;
		12'd3894: data = 1'd0;
		12'd3895: data = 1'd1;
		12'd3896: data = 1'd0;
		12'd3897: data = 1'd1;
		12'd3898: data = 1'd1;
		12'd3899: data = 1'd0;
		12'd3900: data = 1'd1;
		12'd3901: data = 1'd0;
		12'd3902: data = 1'd1;
		12'd3903: data = 1'd0;
		12'd3904: data = 1'd0;
		12'd3905: data = 1'd1;
		12'd3906: data = 1'd1;
		12'd3907: data = 1'd0;
		12'd3908: data = 1'd1;
		12'd3909: data = 1'd0;
		12'd3910: data = 1'd1;
		12'd3911: data = 1'd0;
		12'd3912: data = 1'd1;
		12'd3913: data = 1'd0;
		12'd3914: data = 1'd1;
		12'd3915: data = 1'd0;
		12'd3916: data = 1'd1;
		12'd3917: data = 1'd0;
		12'd3918: data = 1'd1;
		12'd3919: data = 1'd0;
		12'd3920: data = 1'd0;
		12'd3921: data = 1'd1;
		12'd3922: data = 1'd1;
		12'd3923: data = 1'd0;
		12'd3924: data = 1'd1;
		12'd3925: data = 1'd0;
		12'd3926: data = 1'd1;
		12'd3927: data = 1'd0;
		12'd3928: data = 1'd1;
		12'd3929: data = 1'd0;
		12'd3930: data = 1'd1;
		12'd3931: data = 1'd1;
		12'd3932: data = 1'd0;
		12'd3933: data = 1'd1;
		12'd3934: data = 1'd0;
		12'd3935: data = 1'd1;
		12'd3936: data = 1'd0;
		12'd3937: data = 1'd0;
		12'd3938: data = 1'd1;
		12'd3939: data = 1'd1;
		12'd3940: data = 1'd1;
		12'd3941: data = 1'd0;
		12'd3942: data = 1'd1;
		12'd3943: data = 1'd1;
		12'd3944: data = 1'd0;
		12'd3945: data = 1'd1;
		12'd3946: data = 1'd0;
		12'd3947: data = 1'd1;
		12'd3948: data = 1'd0;
		12'd3949: data = 1'd1;
		12'd3950: data = 1'd0;
		12'd3951: data = 1'd1;
		12'd3952: data = 1'd1;
		12'd3953: data = 1'd0;
		12'd3954: data = 1'd1;
		12'd3955: data = 1'd1;
		12'd3956: data = 1'd0;
		12'd3957: data = 1'd1;
		12'd3958: data = 1'd0;
		12'd3959: data = 1'd1;
		12'd3960: data = 1'd0;
		12'd3961: data = 1'd1;
		12'd3962: data = 1'd0;
		12'd3963: data = 1'd1;
		12'd3964: data = 1'd0;
		12'd3965: data = 1'd0;
		12'd3966: data = 1'd1;
		12'd3967: data = 1'd0;
		12'd3968: data = 1'd1;
		12'd3969: data = 1'd0;
		12'd3970: data = 1'd0;
		12'd3971: data = 1'd1;
		12'd3972: data = 1'd0;
		12'd3973: data = 1'd1;
		12'd3974: data = 1'd0;
		12'd3975: data = 1'd1;
		12'd3976: data = 1'd0;
		12'd3977: data = 1'd0;
		12'd3978: data = 1'd1;
		12'd3979: data = 1'd0;
		12'd3980: data = 1'd1;
		12'd3981: data = 1'd0;
		12'd3982: data = 1'd1;
		12'd3983: data = 1'd0;
		12'd3984: data = 1'd1;
		12'd3985: data = 1'd1;
		12'd3986: data = 1'd0;
		12'd3987: data = 1'd1;
		12'd3988: data = 1'd1;
		12'd3989: data = 1'd0;
		12'd3990: data = 1'd1;
		12'd3991: data = 1'd0;
		12'd3992: data = 1'd1;
		12'd3993: data = 1'd0;
		12'd3994: data = 1'd1;
		12'd3995: data = 1'd0;
		12'd3996: data = 1'd1;
		12'd3997: data = 1'd0;
		12'd3998: data = 1'd0;
		12'd3999: data = 1'd1;
		12'd4000: data = 1'd1;
		12'd4001: data = 1'd1;
		12'd4002: data = 1'd0;
		12'd4003: data = 1'd0;
		12'd4004: data = 1'd1;
		12'd4005: data = 1'd0;
		12'd4006: data = 1'd1;
		12'd4007: data = 1'd0;
		12'd4008: data = 1'd1;
		12'd4009: data = 1'd0;
		12'd4010: data = 1'd0;
		12'd4011: data = 1'd1;
		12'd4012: data = 1'd0;
		12'd4013: data = 1'd1;
		12'd4014: data = 1'd0;
		12'd4015: data = 1'd1;
		12'd4016: data = 1'd1;
		12'd4017: data = 1'd1;
		12'd4018: data = 1'd1;
		12'd4019: data = 1'd0;
		12'd4020: data = 1'd1;
		12'd4021: data = 1'd0;
		12'd4022: data = 1'd0;
		12'd4023: data = 1'd1;
		12'd4024: data = 1'd0;
		12'd4025: data = 1'd1;
		12'd4026: data = 1'd0;
		12'd4027: data = 1'd1;
		12'd4028: data = 1'd0;
		12'd4029: data = 1'd1;
		12'd4030: data = 1'd0;
		12'd4031: data = 1'd0;
		12'd4032: data = 1'd1;
		12'd4033: data = 1'd1;
		12'd4034: data = 1'd1;
		12'd4035: data = 1'd0;
		12'd4036: data = 1'd0;
		12'd4037: data = 1'd0;
		12'd4038: data = 1'd0;
		12'd4039: data = 1'd1;
		12'd4040: data = 1'd0;
		12'd4041: data = 1'd1;
		12'd4042: data = 1'd0;
		12'd4043: data = 1'd0;
		12'd4044: data = 1'd1;
		12'd4045: data = 1'd0;
		12'd4046: data = 1'd1;
		12'd4047: data = 1'd0;
		12'd4048: data = 1'd1;
		12'd4049: data = 1'd1;
		12'd4050: data = 1'd1;
		12'd4051: data = 1'd1;
		12'd4052: data = 1'd0;
		12'd4053: data = 1'd0;
		12'd4054: data = 1'd0;
		12'd4055: data = 1'd0;
		12'd4056: data = 1'd1;
		12'd4057: data = 1'd0;
		12'd4058: data = 1'd1;
		12'd4059: data = 1'd0;
		12'd4060: data = 1'd1;
		12'd4061: data = 1'd0;
		12'd4062: data = 1'd1;
		12'd4063: data = 1'd0;
		12'd4064: data = 1'd1;
		12'd4065: data = 1'd1;
		12'd4066: data = 1'd1;
		12'd4067: data = 1'd1;
		12'd4068: data = 1'd0;
		12'd4069: data = 1'd0;
		12'd4070: data = 1'd0;
		12'd4071: data = 1'd0;
		12'd4072: data = 1'd1;
		12'd4073: data = 1'd0;
		12'd4074: data = 1'd1;
		12'd4075: data = 1'd0;
		12'd4076: data = 1'd1;
		12'd4077: data = 1'd0;
		12'd4078: data = 1'd1;
		12'd4079: data = 1'd1;
		12'd4080: data = 1'd1;
		12'd4081: data = 1'd1;
		12'd4082: data = 1'd1;
		12'd4083: data = 1'd1;
		12'd4084: data = 1'd1;
		12'd4085: data = 1'd1;
		12'd4086: data = 1'd1;
		12'd4087: data = 1'd1;
		12'd4088: data = 1'd1;
		12'd4089: data = 1'd0;
		12'd4090: data = 1'd1;
		12'd4091: data = 1'd0;
		12'd4092: data = 1'd0;
		12'd4093: data = 1'd1;
		12'd4094: data = 1'd0;
		12'd4095: data = 1'd1;
		default: data = 1'd0;
	endcase
end
endmodule

module layer0_N7(address, data);
input wire [11:0] address;
output reg [3:0] data;

wire [6:0] i; layer0_N7_idx_1 idx_1_inst(address[11:3], i);
wire [1:0] t; layer0_N7_rsh_1 rsh_1_inst(address[11:3], t);
wire [2:0] b; layer0_N7_2 layer0_N7_2_inst(address[11:3], b);
wire [0:0] lb; layer0_N7_lb_1 lb_1_inst(address, lb);
wire [2:0] u; layer0_N7_ust_1 ust_1_inst({i, address[2:0]}, u);

always @(*) begin
	data = {(u >> t) + b, lb};
end
endmodule
