
module layer1_N0_ust_3(address, data);
input wire [4:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		5'd0: data = 2'd2;
		5'd1: data = 2'd1;
		5'd2: data = 2'd0;
		5'd3: data = 2'd0;
		5'd4: data = 2'd0;
		5'd5: data = 2'd0;
		5'd6: data = 2'd0;
		5'd7: data = 2'd0;
		5'd8: data = 2'd3;
		5'd9: data = 2'd2;
		5'd10: data = 2'd1;
		5'd11: data = 2'd0;
		5'd12: data = 2'd0;
		5'd13: data = 2'd0;
		5'd14: data = 2'd0;
		5'd15: data = 2'd0;
		5'd16: data = 2'd2;
		5'd17: data = 2'd2;
		5'd18: data = 2'd1;
		5'd19: data = 2'd0;
		5'd20: data = 2'd0;
		5'd21: data = 2'd0;
		5'd22: data = 2'd0;
		5'd23: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N0_idx_3(address, data);
input wire [3:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		4'd0: data = 2'd1;
		4'd1: data = 2'd1;
		4'd2: data = 2'd2;
		4'd3: data = 2'd2;
		4'd4: data = 2'd0;
		4'd5: data = 2'd0;
		4'd6: data = 2'd0;
		4'd7: data = 2'd1;
		4'd8: data = 2'd0;
		4'd9: data = 2'd0;
		4'd10: data = 2'd0;
		4'd11: data = 2'd0;
		4'd12: data = 2'd0;
		4'd13: data = 2'd0;
		4'd14: data = 2'd0;
		4'd15: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N0_rsh_3(address, data);
input wire [3:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		4'd0: data = 2'd0;
		4'd1: data = 2'd0;
		4'd2: data = 2'd0;
		4'd3: data = 2'd0;
		4'd4: data = 2'd0;
		4'd5: data = 2'd0;
		4'd6: data = 2'd0;
		4'd7: data = 2'd1;
		4'd8: data = 2'd1;
		4'd9: data = 2'd1;
		4'd10: data = 2'd1;
		4'd11: data = 2'd1;
		4'd12: data = 2'd2;
		4'd13: data = 2'd2;
		4'd14: data = 2'd2;
		4'd15: data = 2'd2;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N0_3(address, data);
input wire [6:0] address;
output reg [1:0] data;

wire [1:0] i; layer1_N0_idx_3 idx_3_inst(address[6:3], i);
wire [1:0] t; layer1_N0_rsh_3 rsh_3_inst(address[6:3], t);
wire [1:0] u; layer1_N0_ust_3 ust_3_inst({i, address[2:0]}, u);

always @(*) begin
	data = (u >> t);
end
endmodule

module layer1_N0_ust_2(address, data);
input wire [7:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		8'd0: data = 2'd3;
		8'd1: data = 2'd2;
		8'd2: data = 2'd1;
		8'd3: data = 2'd0;
		8'd4: data = 2'd3;
		8'd5: data = 2'd2;
		8'd6: data = 2'd1;
		8'd7: data = 2'd0;
		8'd8: data = 2'd2;
		8'd9: data = 2'd1;
		8'd10: data = 2'd0;
		8'd11: data = 2'd0;
		8'd12: data = 2'd2;
		8'd13: data = 2'd1;
		8'd14: data = 2'd0;
		8'd15: data = 2'd0;
		8'd16: data = 2'd2;
		8'd17: data = 2'd1;
		8'd18: data = 2'd1;
		8'd19: data = 2'd0;
		8'd20: data = 2'd2;
		8'd21: data = 2'd1;
		8'd22: data = 2'd0;
		8'd23: data = 2'd0;
		8'd24: data = 2'd2;
		8'd25: data = 2'd1;
		8'd26: data = 2'd1;
		8'd27: data = 2'd1;
		8'd28: data = 2'd2;
		8'd29: data = 2'd1;
		8'd30: data = 2'd1;
		8'd31: data = 2'd0;
		8'd32: data = 2'd3;
		8'd33: data = 2'd3;
		8'd34: data = 2'd2;
		8'd35: data = 2'd0;
		8'd36: data = 2'd3;
		8'd37: data = 2'd3;
		8'd38: data = 2'd2;
		8'd39: data = 2'd0;
		8'd40: data = 2'd3;
		8'd41: data = 2'd2;
		8'd42: data = 2'd1;
		8'd43: data = 2'd1;
		8'd44: data = 2'd3;
		8'd45: data = 2'd2;
		8'd46: data = 2'd1;
		8'd47: data = 2'd0;
		8'd48: data = 2'd3;
		8'd49: data = 2'd2;
		8'd50: data = 2'd0;
		8'd51: data = 2'd0;
		8'd52: data = 2'd3;
		8'd53: data = 2'd1;
		8'd54: data = 2'd0;
		8'd55: data = 2'd0;
		8'd56: data = 2'd2;
		8'd57: data = 2'd0;
		8'd58: data = 2'd0;
		8'd59: data = 2'd0;
		8'd60: data = 2'd2;
		8'd61: data = 2'd0;
		8'd62: data = 2'd0;
		8'd63: data = 2'd0;
		8'd64: data = 2'd2;
		8'd65: data = 2'd1;
		8'd66: data = 2'd1;
		8'd67: data = 2'd0;
		8'd68: data = 2'd2;
		8'd69: data = 2'd1;
		8'd70: data = 2'd1;
		8'd71: data = 2'd0;
		8'd72: data = 2'd2;
		8'd73: data = 2'd0;
		8'd74: data = 2'd0;
		8'd75: data = 2'd0;
		8'd76: data = 2'd2;
		8'd77: data = 2'd1;
		8'd78: data = 2'd0;
		8'd79: data = 2'd0;
		8'd80: data = 2'd2;
		8'd81: data = 2'd2;
		8'd82: data = 2'd1;
		8'd83: data = 2'd1;
		8'd84: data = 2'd2;
		8'd85: data = 2'd2;
		8'd86: data = 2'd1;
		8'd87: data = 2'd0;
		8'd88: data = 2'd3;
		8'd89: data = 2'd2;
		8'd90: data = 2'd2;
		8'd91: data = 2'd1;
		8'd92: data = 2'd3;
		8'd93: data = 2'd2;
		8'd94: data = 2'd1;
		8'd95: data = 2'd0;
		8'd96: data = 2'd3;
		8'd97: data = 2'd2;
		8'd98: data = 2'd2;
		8'd99: data = 2'd0;
		8'd100: data = 2'd3;
		8'd101: data = 2'd3;
		8'd102: data = 2'd2;
		8'd103: data = 2'd0;
		8'd104: data = 2'd3;
		8'd105: data = 2'd2;
		8'd106: data = 2'd1;
		8'd107: data = 2'd0;
		8'd108: data = 2'd3;
		8'd109: data = 2'd3;
		8'd110: data = 2'd2;
		8'd111: data = 2'd0;
		8'd112: data = 2'd3;
		8'd113: data = 2'd1;
		8'd114: data = 2'd0;
		8'd115: data = 2'd0;
		8'd116: data = 2'd3;
		8'd117: data = 2'd1;
		8'd118: data = 2'd0;
		8'd119: data = 2'd0;
		8'd120: data = 2'd2;
		8'd121: data = 2'd1;
		8'd122: data = 2'd1;
		8'd123: data = 2'd0;
		8'd124: data = 2'd3;
		8'd125: data = 2'd2;
		8'd126: data = 2'd1;
		8'd127: data = 2'd0;
		8'd128: data = 2'd2;
		8'd129: data = 2'd1;
		8'd130: data = 2'd0;
		8'd131: data = 2'd0;
		8'd132: data = 2'd2;
		8'd133: data = 2'd0;
		8'd134: data = 2'd0;
		8'd135: data = 2'd0;
		8'd136: data = 2'd2;
		8'd137: data = 2'd0;
		8'd138: data = 2'd0;
		8'd139: data = 2'd0;
		8'd140: data = 2'd1;
		8'd141: data = 2'd0;
		8'd142: data = 2'd0;
		8'd143: data = 2'd0;
		8'd144: data = 2'd3;
		8'd145: data = 2'd2;
		8'd146: data = 2'd1;
		8'd147: data = 2'd0;
		8'd148: data = 2'd3;
		8'd149: data = 2'd2;
		8'd150: data = 2'd2;
		8'd151: data = 2'd0;
		8'd152: data = 2'd1;
		8'd153: data = 2'd1;
		8'd154: data = 2'd1;
		8'd155: data = 2'd1;
		8'd156: data = 2'd1;
		8'd157: data = 2'd1;
		8'd158: data = 2'd0;
		8'd159: data = 2'd1;
		8'd160: data = 2'd2;
		8'd161: data = 2'd2;
		8'd162: data = 2'd1;
		8'd163: data = 2'd0;
		8'd164: data = 2'd2;
		8'd165: data = 2'd2;
		8'd166: data = 2'd1;
		8'd167: data = 2'd0;
		8'd168: data = 2'd1;
		8'd169: data = 2'd1;
		8'd170: data = 2'd1;
		8'd171: data = 2'd1;
		8'd172: data = 2'd1;
		8'd173: data = 2'd1;
		8'd174: data = 2'd0;
		8'd175: data = 2'd0;
		8'd176: data = 2'd1;
		8'd177: data = 2'd1;
		8'd178: data = 2'd0;
		8'd179: data = 2'd1;
		8'd180: data = 2'd1;
		8'd181: data = 2'd1;
		8'd182: data = 2'd0;
		8'd183: data = 2'd0;
		8'd184: data = 2'd3;
		8'd185: data = 2'd2;
		8'd186: data = 2'd1;
		8'd187: data = 2'd0;
		8'd188: data = 2'd3;
		8'd189: data = 2'd2;
		8'd190: data = 2'd0;
		8'd191: data = 2'd0;
		8'd192: data = 2'd3;
		8'd193: data = 2'd2;
		8'd194: data = 2'd0;
		8'd195: data = 2'd0;
		8'd196: data = 2'd3;
		8'd197: data = 2'd2;
		8'd198: data = 2'd0;
		8'd199: data = 2'd0;
		8'd200: data = 2'd3;
		8'd201: data = 2'd1;
		8'd202: data = 2'd0;
		8'd203: data = 2'd0;
		8'd204: data = 2'd3;
		8'd205: data = 2'd2;
		8'd206: data = 2'd1;
		8'd207: data = 2'd0;
		8'd208: data = 2'd3;
		8'd209: data = 2'd1;
		8'd210: data = 2'd0;
		8'd211: data = 2'd0;
		8'd212: data = 2'd3;
		8'd213: data = 2'd1;
		8'd214: data = 2'd1;
		8'd215: data = 2'd0;
		8'd216: data = 2'd2;
		8'd217: data = 2'd1;
		8'd218: data = 2'd0;
		8'd219: data = 2'd0;
		8'd220: data = 2'd3;
		8'd221: data = 2'd1;
		8'd222: data = 2'd0;
		8'd223: data = 2'd0;
		8'd224: data = 2'd2;
		8'd225: data = 2'd1;
		8'd226: data = 2'd0;
		8'd227: data = 2'd0;
		8'd228: data = 2'd2;
		8'd229: data = 2'd1;
		8'd230: data = 2'd1;
		8'd231: data = 2'd0;
		8'd232: data = 2'd2;
		8'd233: data = 2'd1;
		8'd234: data = 2'd0;
		8'd235: data = 2'd0;
		8'd236: data = 2'd2;
		8'd237: data = 2'd2;
		8'd238: data = 2'd1;
		8'd239: data = 2'd0;
		8'd240: data = 2'd1;
		8'd241: data = 2'd0;
		8'd242: data = 2'd0;
		8'd243: data = 2'd0;
		8'd244: data = 2'd2;
		8'd245: data = 2'd0;
		8'd246: data = 2'd0;
		8'd247: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N0_idx_2(address, data);
input wire [6:0] address;
output reg [4:0] data;

always @(*) begin
	case(address)
		7'd0: data = 5'd0;
		7'd1: data = 5'd4;
		7'd2: data = 5'd10;
		7'd3: data = 5'd11;
		7'd4: data = 5'd0;
		7'd5: data = 5'd18;
		7'd6: data = 5'd12;
		7'd7: data = 5'd4;
		7'd8: data = 5'd0;
		7'd9: data = 5'd0;
		7'd10: data = 5'd10;
		7'd11: data = 5'd5;
		7'd12: data = 5'd0;
		7'd13: data = 5'd0;
		7'd14: data = 5'd12;
		7'd15: data = 5'd4;
		7'd16: data = 5'd19;
		7'd17: data = 5'd0;
		7'd18: data = 5'd20;
		7'd19: data = 5'd0;
		7'd20: data = 5'd0;
		7'd21: data = 5'd0;
		7'd22: data = 5'd13;
		7'd23: data = 5'd4;
		7'd24: data = 5'd21;
		7'd25: data = 5'd6;
		7'd26: data = 5'd8;
		7'd27: data = 5'd0;
		7'd28: data = 5'd0;
		7'd29: data = 5'd0;
		7'd30: data = 5'd0;
		7'd31: data = 5'd4;
		7'd32: data = 5'd22;
		7'd33: data = 5'd3;
		7'd34: data = 5'd11;
		7'd35: data = 5'd0;
		7'd36: data = 5'd0;
		7'd37: data = 5'd0;
		7'd38: data = 5'd0;
		7'd39: data = 5'd13;
		7'd40: data = 5'd6;
		7'd41: data = 5'd3;
		7'd42: data = 5'd5;
		7'd43: data = 5'd0;
		7'd44: data = 5'd0;
		7'd45: data = 5'd0;
		7'd46: data = 5'd0;
		7'd47: data = 5'd0;
		7'd48: data = 5'd1;
		7'd49: data = 5'd2;
		7'd50: data = 5'd0;
		7'd51: data = 5'd23;
		7'd52: data = 5'd24;
		7'd53: data = 5'd0;
		7'd54: data = 5'd0;
		7'd55: data = 5'd0;
		7'd56: data = 5'd3;
		7'd57: data = 5'd2;
		7'd58: data = 5'd0;
		7'd59: data = 5'd6;
		7'd60: data = 5'd14;
		7'd61: data = 5'd25;
		7'd62: data = 5'd0;
		7'd63: data = 5'd0;
		7'd64: data = 5'd3;
		7'd65: data = 5'd5;
		7'd66: data = 5'd0;
		7'd67: data = 5'd1;
		7'd68: data = 5'd14;
		7'd69: data = 5'd26;
		7'd70: data = 5'd0;
		7'd71: data = 5'd0;
		7'd72: data = 5'd2;
		7'd73: data = 5'd5;
		7'd74: data = 5'd2;
		7'd75: data = 5'd1;
		7'd76: data = 5'd27;
		7'd77: data = 5'd1;
		7'd78: data = 5'd15;
		7'd79: data = 5'd0;
		7'd80: data = 5'd2;
		7'd81: data = 5'd8;
		7'd82: data = 5'd1;
		7'd83: data = 5'd1;
		7'd84: data = 5'd1;
		7'd85: data = 5'd1;
		7'd86: data = 5'd28;
		7'd87: data = 5'd0;
		7'd88: data = 5'd6;
		7'd89: data = 5'd2;
		7'd90: data = 5'd1;
		7'd91: data = 5'd1;
		7'd92: data = 5'd1;
		7'd93: data = 5'd1;
		7'd94: data = 5'd1;
		7'd95: data = 5'd15;
		7'd96: data = 5'd3;
		7'd97: data = 5'd2;
		7'd98: data = 5'd1;
		7'd99: data = 5'd16;
		7'd100: data = 5'd9;
		7'd101: data = 5'd1;
		7'd102: data = 5'd1;
		7'd103: data = 5'd29;
		7'd104: data = 5'd3;
		7'd105: data = 5'd1;
		7'd106: data = 5'd1;
		7'd107: data = 5'd7;
		7'd108: data = 5'd7;
		7'd109: data = 5'd1;
		7'd110: data = 5'd1;
		7'd111: data = 5'd1;
		7'd112: data = 5'd8;
		7'd113: data = 5'd1;
		7'd114: data = 5'd16;
		7'd115: data = 5'd17;
		7'd116: data = 5'd7;
		7'd117: data = 5'd9;
		7'd118: data = 5'd1;
		7'd119: data = 5'd1;
		7'd120: data = 5'd2;
		7'd121: data = 5'd1;
		7'd122: data = 5'd17;
		7'd123: data = 5'd1;
		7'd124: data = 5'd30;
		7'd125: data = 5'd7;
		7'd126: data = 5'd9;
		7'd127: data = 5'd1;
		default: data = 5'd0;
	endcase
end
endmodule

module layer1_N0_rsh_2(address, data);
input wire [6:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		7'd0: data = 2'd2;
		7'd1: data = 2'd1;
		7'd2: data = 2'd0;
		7'd3: data = 2'd0;
		7'd4: data = 2'd0;
		7'd5: data = 2'd0;
		7'd6: data = 2'd0;
		7'd7: data = 2'd0;
		7'd8: data = 2'd2;
		7'd9: data = 2'd1;
		7'd10: data = 2'd0;
		7'd11: data = 2'd0;
		7'd12: data = 2'd0;
		7'd13: data = 2'd0;
		7'd14: data = 2'd0;
		7'd15: data = 2'd0;
		7'd16: data = 2'd0;
		7'd17: data = 2'd1;
		7'd18: data = 2'd0;
		7'd19: data = 2'd0;
		7'd20: data = 2'd0;
		7'd21: data = 2'd0;
		7'd22: data = 2'd0;
		7'd23: data = 2'd0;
		7'd24: data = 2'd0;
		7'd25: data = 2'd1;
		7'd26: data = 2'd0;
		7'd27: data = 2'd0;
		7'd28: data = 2'd0;
		7'd29: data = 2'd0;
		7'd30: data = 2'd0;
		7'd31: data = 2'd0;
		7'd32: data = 2'd0;
		7'd33: data = 2'd0;
		7'd34: data = 2'd0;
		7'd35: data = 2'd0;
		7'd36: data = 2'd0;
		7'd37: data = 2'd0;
		7'd38: data = 2'd0;
		7'd39: data = 2'd0;
		7'd40: data = 2'd1;
		7'd41: data = 2'd0;
		7'd42: data = 2'd0;
		7'd43: data = 2'd0;
		7'd44: data = 2'd0;
		7'd45: data = 2'd0;
		7'd46: data = 2'd0;
		7'd47: data = 2'd0;
		7'd48: data = 2'd1;
		7'd49: data = 2'd0;
		7'd50: data = 2'd0;
		7'd51: data = 2'd0;
		7'd52: data = 2'd0;
		7'd53: data = 2'd0;
		7'd54: data = 2'd0;
		7'd55: data = 2'd0;
		7'd56: data = 2'd0;
		7'd57: data = 2'd0;
		7'd58: data = 2'd0;
		7'd59: data = 2'd0;
		7'd60: data = 2'd0;
		7'd61: data = 2'd0;
		7'd62: data = 2'd0;
		7'd63: data = 2'd0;
		7'd64: data = 2'd0;
		7'd65: data = 2'd0;
		7'd66: data = 2'd0;
		7'd67: data = 2'd0;
		7'd68: data = 2'd0;
		7'd69: data = 2'd0;
		7'd70: data = 2'd0;
		7'd71: data = 2'd0;
		7'd72: data = 2'd0;
		7'd73: data = 2'd0;
		7'd74: data = 2'd0;
		7'd75: data = 2'd0;
		7'd76: data = 2'd0;
		7'd77: data = 2'd0;
		7'd78: data = 2'd0;
		7'd79: data = 2'd0;
		7'd80: data = 2'd0;
		7'd81: data = 2'd0;
		7'd82: data = 2'd0;
		7'd83: data = 2'd0;
		7'd84: data = 2'd0;
		7'd85: data = 2'd0;
		7'd86: data = 2'd0;
		7'd87: data = 2'd0;
		7'd88: data = 2'd1;
		7'd89: data = 2'd0;
		7'd90: data = 2'd0;
		7'd91: data = 2'd0;
		7'd92: data = 2'd0;
		7'd93: data = 2'd0;
		7'd94: data = 2'd0;
		7'd95: data = 2'd0;
		7'd96: data = 2'd0;
		7'd97: data = 2'd0;
		7'd98: data = 2'd0;
		7'd99: data = 2'd0;
		7'd100: data = 2'd0;
		7'd101: data = 2'd0;
		7'd102: data = 2'd0;
		7'd103: data = 2'd0;
		7'd104: data = 2'd0;
		7'd105: data = 2'd0;
		7'd106: data = 2'd0;
		7'd107: data = 2'd0;
		7'd108: data = 2'd0;
		7'd109: data = 2'd0;
		7'd110: data = 2'd0;
		7'd111: data = 2'd0;
		7'd112: data = 2'd0;
		7'd113: data = 2'd0;
		7'd114: data = 2'd0;
		7'd115: data = 2'd0;
		7'd116: data = 2'd0;
		7'd117: data = 2'd0;
		7'd118: data = 2'd0;
		7'd119: data = 2'd0;
		7'd120: data = 2'd0;
		7'd121: data = 2'd0;
		7'd122: data = 2'd0;
		7'd123: data = 2'd1;
		7'd124: data = 2'd0;
		7'd125: data = 2'd0;
		7'd126: data = 2'd0;
		7'd127: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N0_lb_2(address, data);
input wire [9:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		10'd0: data = 2'd3;
		10'd1: data = 2'd3;
		10'd2: data = 2'd2;
		10'd3: data = 2'd1;
		10'd4: data = 2'd3;
		10'd5: data = 2'd3;
		10'd6: data = 2'd2;
		10'd7: data = 2'd0;
		10'd8: data = 2'd3;
		10'd9: data = 2'd2;
		10'd10: data = 2'd1;
		10'd11: data = 2'd3;
		10'd12: data = 2'd3;
		10'd13: data = 2'd2;
		10'd14: data = 2'd0;
		10'd15: data = 2'd2;
		10'd16: data = 2'd3;
		10'd17: data = 2'd1;
		10'd18: data = 2'd3;
		10'd19: data = 2'd0;
		10'd20: data = 2'd3;
		10'd21: data = 2'd0;
		10'd22: data = 2'd1;
		10'd23: data = 2'd2;
		10'd24: data = 2'd3;
		10'd25: data = 2'd3;
		10'd26: data = 2'd0;
		10'd27: data = 2'd1;
		10'd28: data = 2'd2;
		10'd29: data = 2'd2;
		10'd30: data = 2'd3;
		10'd31: data = 2'd3;
		10'd32: data = 2'd1;
		10'd33: data = 2'd2;
		10'd34: data = 2'd2;
		10'd35: data = 2'd3;
		10'd36: data = 2'd0;
		10'd37: data = 2'd1;
		10'd38: data = 2'd3;
		10'd39: data = 2'd2;
		10'd40: data = 2'd1;
		10'd41: data = 2'd2;
		10'd42: data = 2'd3;
		10'd43: data = 2'd2;
		10'd44: data = 2'd1;
		10'd45: data = 2'd3;
		10'd46: data = 2'd0;
		10'd47: data = 2'd3;
		10'd48: data = 2'd2;
		10'd49: data = 2'd3;
		10'd50: data = 2'd0;
		10'd51: data = 2'd3;
		10'd52: data = 2'd3;
		10'd53: data = 2'd0;
		10'd54: data = 2'd0;
		10'd55: data = 2'd3;
		10'd56: data = 2'd3;
		10'd57: data = 2'd0;
		10'd58: data = 2'd0;
		10'd59: data = 2'd3;
		10'd60: data = 2'd3;
		10'd61: data = 2'd1;
		10'd62: data = 2'd1;
		10'd63: data = 2'd3;
		10'd64: data = 2'd3;
		10'd65: data = 2'd3;
		10'd66: data = 2'd1;
		10'd67: data = 2'd1;
		10'd68: data = 2'd3;
		10'd69: data = 2'd2;
		10'd70: data = 2'd0;
		10'd71: data = 2'd0;
		10'd72: data = 2'd3;
		10'd73: data = 2'd1;
		10'd74: data = 2'd3;
		10'd75: data = 2'd3;
		10'd76: data = 2'd3;
		10'd77: data = 2'd1;
		10'd78: data = 2'd3;
		10'd79: data = 2'd1;
		10'd80: data = 2'd3;
		10'd81: data = 2'd1;
		10'd82: data = 2'd2;
		10'd83: data = 2'd0;
		10'd84: data = 2'd3;
		10'd85: data = 2'd0;
		10'd86: data = 2'd1;
		10'd87: data = 2'd2;
		10'd88: data = 2'd3;
		10'd89: data = 2'd3;
		10'd90: data = 2'd3;
		10'd91: data = 2'd0;
		10'd92: data = 2'd1;
		10'd93: data = 2'd2;
		10'd94: data = 2'd2;
		10'd95: data = 2'd3;
		10'd96: data = 2'd1;
		10'd97: data = 2'd1;
		10'd98: data = 2'd2;
		10'd99: data = 2'd2;
		10'd100: data = 2'd0;
		10'd101: data = 2'd1;
		10'd102: data = 2'd2;
		10'd103: data = 2'd2;
		10'd104: data = 2'd1;
		10'd105: data = 2'd2;
		10'd106: data = 2'd3;
		10'd107: data = 2'd2;
		10'd108: data = 2'd1;
		10'd109: data = 2'd3;
		10'd110: data = 2'd3;
		10'd111: data = 2'd2;
		10'd112: data = 2'd2;
		10'd113: data = 2'd3;
		10'd114: data = 2'd0;
		10'd115: data = 2'd2;
		10'd116: data = 2'd3;
		10'd117: data = 2'd0;
		10'd118: data = 2'd0;
		10'd119: data = 2'd3;
		10'd120: data = 2'd3;
		10'd121: data = 2'd1;
		10'd122: data = 2'd0;
		10'd123: data = 2'd3;
		10'd124: data = 2'd3;
		10'd125: data = 2'd1;
		10'd126: data = 2'd1;
		10'd127: data = 2'd3;
		10'd128: data = 2'd3;
		10'd129: data = 2'd2;
		10'd130: data = 2'd0;
		10'd131: data = 2'd1;
		10'd132: data = 2'd3;
		10'd133: data = 2'd1;
		10'd134: data = 2'd3;
		10'd135: data = 2'd0;
		10'd136: data = 2'd3;
		10'd137: data = 2'd1;
		10'd138: data = 2'd2;
		10'd139: data = 2'd2;
		10'd140: data = 2'd3;
		10'd141: data = 2'd0;
		10'd142: data = 2'd2;
		10'd143: data = 2'd0;
		10'd144: data = 2'd3;
		10'd145: data = 2'd0;
		10'd146: data = 2'd1;
		10'd147: data = 2'd3;
		10'd148: data = 2'd3;
		10'd149: data = 2'd0;
		10'd150: data = 2'd1;
		10'd151: data = 2'd1;
		10'd152: data = 2'd2;
		10'd153: data = 2'd3;
		10'd154: data = 2'd3;
		10'd155: data = 2'd3;
		10'd156: data = 2'd1;
		10'd157: data = 2'd2;
		10'd158: data = 2'd2;
		10'd159: data = 2'd2;
		10'd160: data = 2'd0;
		10'd161: data = 2'd1;
		10'd162: data = 2'd1;
		10'd163: data = 2'd1;
		10'd164: data = 2'd0;
		10'd165: data = 2'd1;
		10'd166: data = 2'd2;
		10'd167: data = 2'd1;
		10'd168: data = 2'd1;
		10'd169: data = 2'd2;
		10'd170: data = 2'd2;
		10'd171: data = 2'd2;
		10'd172: data = 2'd1;
		10'd173: data = 2'd2;
		10'd174: data = 2'd3;
		10'd175: data = 2'd2;
		10'd176: data = 2'd2;
		10'd177: data = 2'd3;
		10'd178: data = 2'd3;
		10'd179: data = 2'd2;
		10'd180: data = 2'd3;
		10'd181: data = 2'd0;
		10'd182: data = 2'd0;
		10'd183: data = 2'd2;
		10'd184: data = 2'd3;
		10'd185: data = 2'd0;
		10'd186: data = 2'd0;
		10'd187: data = 2'd3;
		10'd188: data = 2'd3;
		10'd189: data = 2'd1;
		10'd190: data = 2'd1;
		10'd191: data = 2'd3;
		10'd192: data = 2'd3;
		10'd193: data = 2'd1;
		10'd194: data = 2'd0;
		10'd195: data = 2'd0;
		10'd196: data = 2'd3;
		10'd197: data = 2'd1;
		10'd198: data = 2'd3;
		10'd199: data = 2'd3;
		10'd200: data = 2'd3;
		10'd201: data = 2'd0;
		10'd202: data = 2'd2;
		10'd203: data = 2'd1;
		10'd204: data = 2'd3;
		10'd205: data = 2'd3;
		10'd206: data = 2'd1;
		10'd207: data = 2'd0;
		10'd208: data = 2'd3;
		10'd209: data = 2'd3;
		10'd210: data = 2'd1;
		10'd211: data = 2'd2;
		10'd212: data = 2'd3;
		10'd213: data = 2'd3;
		10'd214: data = 2'd0;
		10'd215: data = 2'd0;
		10'd216: data = 2'd2;
		10'd217: data = 2'd2;
		10'd218: data = 2'd3;
		10'd219: data = 2'd2;
		10'd220: data = 2'd1;
		10'd221: data = 2'd1;
		10'd222: data = 2'd1;
		10'd223: data = 2'd1;
		10'd224: data = 2'd0;
		10'd225: data = 2'd1;
		10'd226: data = 2'd1;
		10'd227: data = 2'd1;
		10'd228: data = 2'd0;
		10'd229: data = 2'd1;
		10'd230: data = 2'd1;
		10'd231: data = 2'd0;
		10'd232: data = 2'd1;
		10'd233: data = 2'd1;
		10'd234: data = 2'd2;
		10'd235: data = 2'd1;
		10'd236: data = 2'd1;
		10'd237: data = 2'd2;
		10'd238: data = 2'd2;
		10'd239: data = 2'd2;
		10'd240: data = 2'd2;
		10'd241: data = 2'd2;
		10'd242: data = 2'd3;
		10'd243: data = 2'd2;
		10'd244: data = 2'd2;
		10'd245: data = 2'd3;
		10'd246: data = 2'd3;
		10'd247: data = 2'd2;
		10'd248: data = 2'd3;
		10'd249: data = 2'd0;
		10'd250: data = 2'd0;
		10'd251: data = 2'd2;
		10'd252: data = 2'd3;
		10'd253: data = 2'd0;
		10'd254: data = 2'd0;
		10'd255: data = 2'd3;
		10'd256: data = 2'd3;
		10'd257: data = 2'd0;
		10'd258: data = 2'd3;
		10'd259: data = 2'd0;
		10'd260: data = 2'd3;
		10'd261: data = 2'd0;
		10'd262: data = 2'd2;
		10'd263: data = 2'd2;
		10'd264: data = 2'd3;
		10'd265: data = 2'd3;
		10'd266: data = 2'd1;
		10'd267: data = 2'd0;
		10'd268: data = 2'd3;
		10'd269: data = 2'd3;
		10'd270: data = 2'd1;
		10'd271: data = 2'd3;
		10'd272: data = 2'd2;
		10'd273: data = 2'd2;
		10'd274: data = 2'd0;
		10'd275: data = 2'd1;
		10'd276: data = 2'd2;
		10'd277: data = 2'd2;
		10'd278: data = 2'd3;
		10'd279: data = 2'd3;
		10'd280: data = 2'd2;
		10'd281: data = 2'd2;
		10'd282: data = 2'd2;
		10'd283: data = 2'd2;
		10'd284: data = 2'd1;
		10'd285: data = 2'd1;
		10'd286: data = 2'd1;
		10'd287: data = 2'd1;
		10'd288: data = 2'd0;
		10'd289: data = 2'd0;
		10'd290: data = 2'd1;
		10'd291: data = 2'd0;
		10'd292: data = 2'd0;
		10'd293: data = 2'd0;
		10'd294: data = 2'd1;
		10'd295: data = 2'd0;
		10'd296: data = 2'd0;
		10'd297: data = 2'd1;
		10'd298: data = 2'd1;
		10'd299: data = 2'd0;
		10'd300: data = 2'd1;
		10'd301: data = 2'd1;
		10'd302: data = 2'd2;
		10'd303: data = 2'd1;
		10'd304: data = 2'd1;
		10'd305: data = 2'd2;
		10'd306: data = 2'd2;
		10'd307: data = 2'd2;
		10'd308: data = 2'd2;
		10'd309: data = 2'd3;
		10'd310: data = 2'd3;
		10'd311: data = 2'd2;
		10'd312: data = 2'd3;
		10'd313: data = 2'd3;
		10'd314: data = 2'd3;
		10'd315: data = 2'd2;
		10'd316: data = 2'd3;
		10'd317: data = 2'd0;
		10'd318: data = 2'd0;
		10'd319: data = 2'd3;
		10'd320: data = 2'd3;
		10'd321: data = 2'd0;
		10'd322: data = 2'd3;
		10'd323: data = 2'd3;
		10'd324: data = 2'd3;
		10'd325: data = 2'd3;
		10'd326: data = 2'd2;
		10'd327: data = 2'd1;
		10'd328: data = 2'd2;
		10'd329: data = 2'd3;
		10'd330: data = 2'd1;
		10'd331: data = 2'd0;
		10'd332: data = 2'd2;
		10'd333: data = 2'd2;
		10'd334: data = 2'd0;
		10'd335: data = 2'd2;
		10'd336: data = 2'd2;
		10'd337: data = 2'd2;
		10'd338: data = 2'd3;
		10'd339: data = 2'd0;
		10'd340: data = 2'd1;
		10'd341: data = 2'd2;
		10'd342: data = 2'd2;
		10'd343: data = 2'd2;
		10'd344: data = 2'd1;
		10'd345: data = 2'd1;
		10'd346: data = 2'd1;
		10'd347: data = 2'd1;
		10'd348: data = 2'd1;
		10'd349: data = 2'd1;
		10'd350: data = 2'd0;
		10'd351: data = 2'd0;
		10'd352: data = 2'd0;
		10'd353: data = 2'd0;
		10'd354: data = 2'd0;
		10'd355: data = 2'd0;
		10'd356: data = 2'd0;
		10'd357: data = 2'd0;
		10'd358: data = 2'd0;
		10'd359: data = 2'd0;
		10'd360: data = 2'd0;
		10'd361: data = 2'd0;
		10'd362: data = 2'd1;
		10'd363: data = 2'd0;
		10'd364: data = 2'd0;
		10'd365: data = 2'd1;
		10'd366: data = 2'd1;
		10'd367: data = 2'd1;
		10'd368: data = 2'd1;
		10'd369: data = 2'd1;
		10'd370: data = 2'd2;
		10'd371: data = 2'd1;
		10'd372: data = 2'd2;
		10'd373: data = 2'd2;
		10'd374: data = 2'd2;
		10'd375: data = 2'd2;
		10'd376: data = 2'd2;
		10'd377: data = 2'd3;
		10'd378: data = 2'd3;
		10'd379: data = 2'd2;
		10'd380: data = 2'd3;
		10'd381: data = 2'd3;
		10'd382: data = 2'd3;
		10'd383: data = 2'd3;
		10'd384: data = 2'd2;
		10'd385: data = 2'd3;
		10'd386: data = 2'd2;
		10'd387: data = 2'd2;
		10'd388: data = 2'd2;
		10'd389: data = 2'd2;
		10'd390: data = 2'd1;
		10'd391: data = 2'd0;
		10'd392: data = 2'd2;
		10'd393: data = 2'd2;
		10'd394: data = 2'd0;
		10'd395: data = 2'd3;
		10'd396: data = 2'd2;
		10'd397: data = 2'd1;
		10'd398: data = 2'd3;
		10'd399: data = 2'd1;
		10'd400: data = 2'd1;
		10'd401: data = 2'd1;
		10'd402: data = 2'd3;
		10'd403: data = 2'd3;
		10'd404: data = 2'd1;
		10'd405: data = 2'd1;
		10'd406: data = 2'd2;
		10'd407: data = 2'd1;
		10'd408: data = 2'd1;
		10'd409: data = 2'd1;
		10'd410: data = 2'd0;
		10'd411: data = 2'd1;
		10'd412: data = 2'd0;
		10'd413: data = 2'd0;
		10'd414: data = 2'd3;
		10'd415: data = 2'd0;
		10'd416: data = 2'd0;
		10'd417: data = 2'd0;
		10'd418: data = 2'd3;
		10'd419: data = 2'd0;
		10'd420: data = 2'd0;
		10'd421: data = 2'd0;
		10'd422: data = 2'd3;
		10'd423: data = 2'd0;
		10'd424: data = 2'd0;
		10'd425: data = 2'd0;
		10'd426: data = 2'd0;
		10'd427: data = 2'd0;
		10'd428: data = 2'd0;
		10'd429: data = 2'd0;
		10'd430: data = 2'd1;
		10'd431: data = 2'd0;
		10'd432: data = 2'd1;
		10'd433: data = 2'd1;
		10'd434: data = 2'd1;
		10'd435: data = 2'd1;
		10'd436: data = 2'd1;
		10'd437: data = 2'd1;
		10'd438: data = 2'd2;
		10'd439: data = 2'd1;
		10'd440: data = 2'd2;
		10'd441: data = 2'd2;
		10'd442: data = 2'd2;
		10'd443: data = 2'd2;
		10'd444: data = 2'd2;
		10'd445: data = 2'd3;
		10'd446: data = 2'd3;
		10'd447: data = 2'd2;
		10'd448: data = 2'd2;
		10'd449: data = 2'd2;
		10'd450: data = 2'd2;
		10'd451: data = 2'd1;
		10'd452: data = 2'd2;
		10'd453: data = 2'd2;
		10'd454: data = 2'd1;
		10'd455: data = 2'd3;
		10'd456: data = 2'd1;
		10'd457: data = 2'd1;
		10'd458: data = 2'd0;
		10'd459: data = 2'd2;
		10'd460: data = 2'd1;
		10'd461: data = 2'd1;
		10'd462: data = 2'd3;
		10'd463: data = 2'd0;
		10'd464: data = 2'd1;
		10'd465: data = 2'd1;
		10'd466: data = 2'd2;
		10'd467: data = 2'd2;
		10'd468: data = 2'd0;
		10'd469: data = 2'd0;
		10'd470: data = 2'd1;
		10'd471: data = 2'd1;
		10'd472: data = 2'd0;
		10'd473: data = 2'd0;
		10'd474: data = 2'd3;
		10'd475: data = 2'd0;
		10'd476: data = 2'd0;
		10'd477: data = 2'd3;
		10'd478: data = 2'd2;
		10'd479: data = 2'd0;
		10'd480: data = 2'd0;
		10'd481: data = 2'd3;
		10'd482: data = 2'd2;
		10'd483: data = 2'd0;
		10'd484: data = 2'd0;
		10'd485: data = 2'd3;
		10'd486: data = 2'd2;
		10'd487: data = 2'd0;
		10'd488: data = 2'd0;
		10'd489: data = 2'd3;
		10'd490: data = 2'd3;
		10'd491: data = 2'd0;
		10'd492: data = 2'd0;
		10'd493: data = 2'd0;
		10'd494: data = 2'd0;
		10'd495: data = 2'd0;
		10'd496: data = 2'd0;
		10'd497: data = 2'd0;
		10'd498: data = 2'd1;
		10'd499: data = 2'd0;
		10'd500: data = 2'd1;
		10'd501: data = 2'd1;
		10'd502: data = 2'd1;
		10'd503: data = 2'd1;
		10'd504: data = 2'd1;
		10'd505: data = 2'd2;
		10'd506: data = 2'd2;
		10'd507: data = 2'd1;
		10'd508: data = 2'd2;
		10'd509: data = 2'd2;
		10'd510: data = 2'd3;
		10'd511: data = 2'd2;
		10'd512: data = 2'd1;
		10'd513: data = 2'd2;
		10'd514: data = 2'd1;
		10'd515: data = 2'd0;
		10'd516: data = 2'd1;
		10'd517: data = 2'd1;
		10'd518: data = 2'd0;
		10'd519: data = 2'd3;
		10'd520: data = 2'd1;
		10'd521: data = 2'd1;
		10'd522: data = 2'd3;
		10'd523: data = 2'd1;
		10'd524: data = 2'd0;
		10'd525: data = 2'd0;
		10'd526: data = 2'd2;
		10'd527: data = 2'd3;
		10'd528: data = 2'd0;
		10'd529: data = 2'd0;
		10'd530: data = 2'd1;
		10'd531: data = 2'd2;
		10'd532: data = 2'd0;
		10'd533: data = 2'd0;
		10'd534: data = 2'd0;
		10'd535: data = 2'd0;
		10'd536: data = 2'd3;
		10'd537: data = 2'd3;
		10'd538: data = 2'd2;
		10'd539: data = 2'd0;
		10'd540: data = 2'd3;
		10'd541: data = 2'd2;
		10'd542: data = 2'd1;
		10'd543: data = 2'd0;
		10'd544: data = 2'd0;
		10'd545: data = 2'd2;
		10'd546: data = 2'd1;
		10'd547: data = 2'd0;
		10'd548: data = 2'd0;
		10'd549: data = 2'd3;
		10'd550: data = 2'd2;
		10'd551: data = 2'd0;
		10'd552: data = 2'd0;
		10'd553: data = 2'd3;
		10'd554: data = 2'd2;
		10'd555: data = 2'd0;
		10'd556: data = 2'd0;
		10'd557: data = 2'd3;
		10'd558: data = 2'd0;
		10'd559: data = 2'd0;
		10'd560: data = 2'd0;
		10'd561: data = 2'd0;
		10'd562: data = 2'd0;
		10'd563: data = 2'd0;
		10'd564: data = 2'd0;
		10'd565: data = 2'd0;
		10'd566: data = 2'd1;
		10'd567: data = 2'd0;
		10'd568: data = 2'd1;
		10'd569: data = 2'd1;
		10'd570: data = 2'd1;
		10'd571: data = 2'd1;
		10'd572: data = 2'd2;
		10'd573: data = 2'd2;
		10'd574: data = 2'd2;
		10'd575: data = 2'd1;
		10'd576: data = 2'd1;
		10'd577: data = 2'd1;
		10'd578: data = 2'd1;
		10'd579: data = 2'd3;
		10'd580: data = 2'd0;
		10'd581: data = 2'd1;
		10'd582: data = 2'd3;
		10'd583: data = 2'd2;
		10'd584: data = 2'd0;
		10'd585: data = 2'd0;
		10'd586: data = 2'd2;
		10'd587: data = 2'd0;
		10'd588: data = 2'd0;
		10'd589: data = 2'd0;
		10'd590: data = 2'd1;
		10'd591: data = 2'd2;
		10'd592: data = 2'd3;
		10'd593: data = 2'd3;
		10'd594: data = 2'd0;
		10'd595: data = 2'd1;
		10'd596: data = 2'd3;
		10'd597: data = 2'd3;
		10'd598: data = 2'd3;
		10'd599: data = 2'd0;
		10'd600: data = 2'd3;
		10'd601: data = 2'd2;
		10'd602: data = 2'd2;
		10'd603: data = 2'd0;
		10'd604: data = 2'd3;
		10'd605: data = 2'd2;
		10'd606: data = 2'd1;
		10'd607: data = 2'd0;
		10'd608: data = 2'd3;
		10'd609: data = 2'd2;
		10'd610: data = 2'd1;
		10'd611: data = 2'd0;
		10'd612: data = 2'd0;
		10'd613: data = 2'd2;
		10'd614: data = 2'd1;
		10'd615: data = 2'd0;
		10'd616: data = 2'd3;
		10'd617: data = 2'd3;
		10'd618: data = 2'd2;
		10'd619: data = 2'd0;
		10'd620: data = 2'd3;
		10'd621: data = 2'd3;
		10'd622: data = 2'd3;
		10'd623: data = 2'd0;
		10'd624: data = 2'd3;
		10'd625: data = 2'd3;
		10'd626: data = 2'd0;
		10'd627: data = 2'd0;
		10'd628: data = 2'd0;
		10'd629: data = 2'd0;
		10'd630: data = 2'd0;
		10'd631: data = 2'd0;
		10'd632: data = 2'd0;
		10'd633: data = 2'd0;
		10'd634: data = 2'd1;
		10'd635: data = 2'd0;
		10'd636: data = 2'd1;
		10'd637: data = 2'd1;
		10'd638: data = 2'd2;
		10'd639: data = 2'd1;
		10'd640: data = 2'd0;
		10'd641: data = 2'd0;
		10'd642: data = 2'd0;
		10'd643: data = 2'd3;
		10'd644: data = 2'd0;
		10'd645: data = 2'd0;
		10'd646: data = 2'd3;
		10'd647: data = 2'd1;
		10'd648: data = 2'd3;
		10'd649: data = 2'd3;
		10'd650: data = 2'd1;
		10'd651: data = 2'd3;
		10'd652: data = 2'd3;
		10'd653: data = 2'd3;
		10'd654: data = 2'd0;
		10'd655: data = 2'd2;
		10'd656: data = 2'd3;
		10'd657: data = 2'd3;
		10'd658: data = 2'd3;
		10'd659: data = 2'd0;
		10'd660: data = 2'd2;
		10'd661: data = 2'd2;
		10'd662: data = 2'd2;
		10'd663: data = 2'd0;
		10'd664: data = 2'd2;
		10'd665: data = 2'd1;
		10'd666: data = 2'd1;
		10'd667: data = 2'd0;
		10'd668: data = 2'd2;
		10'd669: data = 2'd1;
		10'd670: data = 2'd0;
		10'd671: data = 2'd0;
		10'd672: data = 2'd3;
		10'd673: data = 2'd1;
		10'd674: data = 2'd0;
		10'd675: data = 2'd0;
		10'd676: data = 2'd3;
		10'd677: data = 2'd1;
		10'd678: data = 2'd0;
		10'd679: data = 2'd0;
		10'd680: data = 2'd3;
		10'd681: data = 2'd2;
		10'd682: data = 2'd1;
		10'd683: data = 2'd0;
		10'd684: data = 2'd3;
		10'd685: data = 2'd3;
		10'd686: data = 2'd2;
		10'd687: data = 2'd0;
		10'd688: data = 2'd3;
		10'd689: data = 2'd3;
		10'd690: data = 2'd3;
		10'd691: data = 2'd0;
		10'd692: data = 2'd3;
		10'd693: data = 2'd3;
		10'd694: data = 2'd0;
		10'd695: data = 2'd0;
		10'd696: data = 2'd0;
		10'd697: data = 2'd0;
		10'd698: data = 2'd0;
		10'd699: data = 2'd0;
		10'd700: data = 2'd1;
		10'd701: data = 2'd1;
		10'd702: data = 2'd1;
		10'd703: data = 2'd1;
		10'd704: data = 2'd3;
		10'd705: data = 2'd0;
		10'd706: data = 2'd3;
		10'd707: data = 2'd2;
		10'd708: data = 2'd3;
		10'd709: data = 2'd3;
		10'd710: data = 2'd2;
		10'd711: data = 2'd0;
		10'd712: data = 2'd3;
		10'd713: data = 2'd3;
		10'd714: data = 2'd1;
		10'd715: data = 2'd2;
		10'd716: data = 2'd2;
		10'd717: data = 2'd2;
		10'd718: data = 2'd3;
		10'd719: data = 2'd1;
		10'd720: data = 2'd2;
		10'd721: data = 2'd2;
		10'd722: data = 2'd2;
		10'd723: data = 2'd0;
		10'd724: data = 2'd2;
		10'd725: data = 2'd1;
		10'd726: data = 2'd1;
		10'd727: data = 2'd0;
		10'd728: data = 2'd2;
		10'd729: data = 2'd1;
		10'd730: data = 2'd0;
		10'd731: data = 2'd0;
		10'd732: data = 2'd2;
		10'd733: data = 2'd0;
		10'd734: data = 2'd0;
		10'd735: data = 2'd0;
		10'd736: data = 2'd2;
		10'd737: data = 2'd0;
		10'd738: data = 2'd0;
		10'd739: data = 2'd0;
		10'd740: data = 2'd3;
		10'd741: data = 2'd1;
		10'd742: data = 2'd0;
		10'd743: data = 2'd0;
		10'd744: data = 2'd3;
		10'd745: data = 2'd1;
		10'd746: data = 2'd0;
		10'd747: data = 2'd0;
		10'd748: data = 2'd3;
		10'd749: data = 2'd2;
		10'd750: data = 2'd1;
		10'd751: data = 2'd0;
		10'd752: data = 2'd3;
		10'd753: data = 2'd2;
		10'd754: data = 2'd2;
		10'd755: data = 2'd0;
		10'd756: data = 2'd3;
		10'd757: data = 2'd3;
		10'd758: data = 2'd3;
		10'd759: data = 2'd0;
		10'd760: data = 2'd3;
		10'd761: data = 2'd3;
		10'd762: data = 2'd0;
		10'd763: data = 2'd0;
		10'd764: data = 2'd0;
		10'd765: data = 2'd0;
		10'd766: data = 2'd1;
		10'd767: data = 2'd0;
		10'd768: data = 2'd3;
		10'd769: data = 2'd3;
		10'd770: data = 2'd3;
		10'd771: data = 2'd1;
		10'd772: data = 2'd2;
		10'd773: data = 2'd3;
		10'd774: data = 2'd1;
		10'd775: data = 2'd3;
		10'd776: data = 2'd2;
		10'd777: data = 2'd2;
		10'd778: data = 2'd0;
		10'd779: data = 2'd2;
		10'd780: data = 2'd2;
		10'd781: data = 2'd2;
		10'd782: data = 2'd2;
		10'd783: data = 2'd1;
		10'd784: data = 2'd1;
		10'd785: data = 2'd1;
		10'd786: data = 2'd1;
		10'd787: data = 2'd0;
		10'd788: data = 2'd1;
		10'd789: data = 2'd1;
		10'd790: data = 2'd0;
		10'd791: data = 2'd0;
		10'd792: data = 2'd1;
		10'd793: data = 2'd0;
		10'd794: data = 2'd0;
		10'd795: data = 2'd0;
		10'd796: data = 2'd1;
		10'd797: data = 2'd3;
		10'd798: data = 2'd0;
		10'd799: data = 2'd0;
		10'd800: data = 2'd1;
		10'd801: data = 2'd3;
		10'd802: data = 2'd0;
		10'd803: data = 2'd0;
		10'd804: data = 2'd2;
		10'd805: data = 2'd0;
		10'd806: data = 2'd0;
		10'd807: data = 2'd0;
		10'd808: data = 2'd3;
		10'd809: data = 2'd1;
		10'd810: data = 2'd0;
		10'd811: data = 2'd0;
		10'd812: data = 2'd3;
		10'd813: data = 2'd1;
		10'd814: data = 2'd0;
		10'd815: data = 2'd0;
		10'd816: data = 2'd3;
		10'd817: data = 2'd2;
		10'd818: data = 2'd1;
		10'd819: data = 2'd0;
		10'd820: data = 2'd3;
		10'd821: data = 2'd2;
		10'd822: data = 2'd2;
		10'd823: data = 2'd0;
		10'd824: data = 2'd3;
		10'd825: data = 2'd3;
		10'd826: data = 2'd3;
		10'd827: data = 2'd0;
		10'd828: data = 2'd3;
		10'd829: data = 2'd0;
		10'd830: data = 2'd0;
		10'd831: data = 2'd0;
		10'd832: data = 2'd2;
		10'd833: data = 2'd3;
		10'd834: data = 2'd2;
		10'd835: data = 2'd0;
		10'd836: data = 2'd2;
		10'd837: data = 2'd2;
		10'd838: data = 2'd0;
		10'd839: data = 2'd3;
		10'd840: data = 2'd1;
		10'd841: data = 2'd1;
		10'd842: data = 2'd3;
		10'd843: data = 2'd1;
		10'd844: data = 2'd1;
		10'd845: data = 2'd1;
		10'd846: data = 2'd1;
		10'd847: data = 2'd0;
		10'd848: data = 2'd1;
		10'd849: data = 2'd1;
		10'd850: data = 2'd0;
		10'd851: data = 2'd0;
		10'd852: data = 2'd1;
		10'd853: data = 2'd0;
		10'd854: data = 2'd0;
		10'd855: data = 2'd0;
		10'd856: data = 2'd0;
		10'd857: data = 2'd3;
		10'd858: data = 2'd0;
		10'd859: data = 2'd0;
		10'd860: data = 2'd0;
		10'd861: data = 2'd2;
		10'd862: data = 2'd0;
		10'd863: data = 2'd0;
		10'd864: data = 2'd0;
		10'd865: data = 2'd2;
		10'd866: data = 2'd0;
		10'd867: data = 2'd0;
		10'd868: data = 2'd1;
		10'd869: data = 2'd3;
		10'd870: data = 2'd0;
		10'd871: data = 2'd0;
		10'd872: data = 2'd2;
		10'd873: data = 2'd0;
		10'd874: data = 2'd0;
		10'd875: data = 2'd0;
		10'd876: data = 2'd2;
		10'd877: data = 2'd0;
		10'd878: data = 2'd0;
		10'd879: data = 2'd0;
		10'd880: data = 2'd2;
		10'd881: data = 2'd1;
		10'd882: data = 2'd0;
		10'd883: data = 2'd0;
		10'd884: data = 2'd2;
		10'd885: data = 2'd2;
		10'd886: data = 2'd1;
		10'd887: data = 2'd0;
		10'd888: data = 2'd2;
		10'd889: data = 2'd3;
		10'd890: data = 2'd2;
		10'd891: data = 2'd0;
		10'd892: data = 2'd3;
		10'd893: data = 2'd3;
		10'd894: data = 2'd3;
		10'd895: data = 2'd0;
		10'd896: data = 2'd1;
		10'd897: data = 2'd2;
		10'd898: data = 2'd1;
		10'd899: data = 2'd3;
		10'd900: data = 2'd1;
		10'd901: data = 2'd1;
		10'd902: data = 2'd0;
		10'd903: data = 2'd2;
		10'd904: data = 2'd1;
		10'd905: data = 2'd1;
		10'd906: data = 2'd2;
		10'd907: data = 2'd1;
		10'd908: data = 2'd0;
		10'd909: data = 2'd0;
		10'd910: data = 2'd0;
		10'd911: data = 2'd0;
		10'd912: data = 2'd0;
		10'd913: data = 2'd0;
		10'd914: data = 2'd0;
		10'd915: data = 2'd0;
		10'd916: data = 2'd0;
		10'd917: data = 2'd3;
		10'd918: data = 2'd0;
		10'd919: data = 2'd0;
		10'd920: data = 2'd0;
		10'd921: data = 2'd2;
		10'd922: data = 2'd0;
		10'd923: data = 2'd0;
		10'd924: data = 2'd3;
		10'd925: data = 2'd1;
		10'd926: data = 2'd0;
		10'd927: data = 2'd0;
		10'd928: data = 2'd0;
		10'd929: data = 2'd2;
		10'd930: data = 2'd0;
		10'd931: data = 2'd0;
		10'd932: data = 2'd0;
		10'd933: data = 2'd2;
		10'd934: data = 2'd0;
		10'd935: data = 2'd0;
		10'd936: data = 2'd1;
		10'd937: data = 2'd3;
		10'd938: data = 2'd0;
		10'd939: data = 2'd0;
		10'd940: data = 2'd2;
		10'd941: data = 2'd0;
		10'd942: data = 2'd0;
		10'd943: data = 2'd0;
		10'd944: data = 2'd2;
		10'd945: data = 2'd0;
		10'd946: data = 2'd0;
		10'd947: data = 2'd0;
		10'd948: data = 2'd2;
		10'd949: data = 2'd1;
		10'd950: data = 2'd0;
		10'd951: data = 2'd0;
		10'd952: data = 2'd2;
		10'd953: data = 2'd2;
		10'd954: data = 2'd1;
		10'd955: data = 2'd0;
		10'd956: data = 2'd2;
		10'd957: data = 2'd3;
		10'd958: data = 2'd2;
		10'd959: data = 2'd0;
		10'd960: data = 2'd1;
		10'd961: data = 2'd1;
		10'd962: data = 2'd0;
		10'd963: data = 2'd3;
		10'd964: data = 2'd0;
		10'd965: data = 2'd1;
		10'd966: data = 2'd3;
		10'd967: data = 2'd1;
		10'd968: data = 2'd0;
		10'd969: data = 2'd0;
		10'd970: data = 2'd1;
		10'd971: data = 2'd0;
		10'd972: data = 2'd0;
		10'd973: data = 2'd0;
		10'd974: data = 2'd0;
		10'd975: data = 2'd0;
		10'd976: data = 2'd0;
		10'd977: data = 2'd3;
		10'd978: data = 2'd0;
		10'd979: data = 2'd0;
		10'd980: data = 2'd3;
		10'd981: data = 2'd2;
		10'd982: data = 2'd0;
		10'd983: data = 2'd0;
		10'd984: data = 2'd3;
		10'd985: data = 2'd1;
		10'd986: data = 2'd0;
		10'd987: data = 2'd0;
		10'd988: data = 2'd2;
		10'd989: data = 2'd0;
		10'd990: data = 2'd0;
		10'd991: data = 2'd0;
		10'd992: data = 2'd3;
		10'd993: data = 2'd1;
		10'd994: data = 2'd0;
		10'd995: data = 2'd0;
		10'd996: data = 2'd0;
		10'd997: data = 2'd2;
		10'd998: data = 2'd0;
		10'd999: data = 2'd0;
		10'd1000: data = 2'd0;
		10'd1001: data = 2'd2;
		10'd1002: data = 2'd0;
		10'd1003: data = 2'd0;
		10'd1004: data = 2'd1;
		10'd1005: data = 2'd3;
		10'd1006: data = 2'd0;
		10'd1007: data = 2'd0;
		10'd1008: data = 2'd1;
		10'd1009: data = 2'd3;
		10'd1010: data = 2'd0;
		10'd1011: data = 2'd0;
		10'd1012: data = 2'd2;
		10'd1013: data = 2'd0;
		10'd1014: data = 2'd0;
		10'd1015: data = 2'd0;
		10'd1016: data = 2'd2;
		10'd1017: data = 2'd1;
		10'd1018: data = 2'd0;
		10'd1019: data = 2'd0;
		10'd1020: data = 2'd2;
		10'd1021: data = 2'd2;
		10'd1022: data = 2'd1;
		10'd1023: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N0_2(address, data);
input wire [9:0] address;
output reg [3:0] data;

wire [4:0] i; layer1_N0_idx_2 idx_2_inst(address[9:3], i);
wire [1:0] t; layer1_N0_rsh_2 rsh_2_inst(address[9:3], t);
wire [1:0] b; layer1_N0_3 layer1_N0_3_inst(address[9:3], b);
wire [1:0] lb; layer1_N0_lb_2 lb_2_inst(address, lb);
wire [1:0] u; layer1_N0_ust_2 ust_2_inst({i, address[2:0]}, u);

always @(*) begin
	data = {(u >> t) + b, lb};
end
endmodule

module layer1_N0_ust_1(address, data);
input wire [6:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		7'd0: data = 3'd6;
		7'd1: data = 3'd4;
		7'd2: data = 3'd2;
		7'd3: data = 3'd0;
		7'd4: data = 3'd4;
		7'd5: data = 3'd3;
		7'd6: data = 3'd1;
		7'd7: data = 3'd0;
		7'd8: data = 3'd4;
		7'd9: data = 3'd3;
		7'd10: data = 3'd2;
		7'd11: data = 3'd0;
		7'd12: data = 3'd5;
		7'd13: data = 3'd4;
		7'd14: data = 3'd2;
		7'd15: data = 3'd0;
		7'd16: data = 3'd4;
		7'd17: data = 3'd2;
		7'd18: data = 3'd1;
		7'd19: data = 3'd0;
		7'd20: data = 3'd3;
		7'd21: data = 3'd3;
		7'd22: data = 3'd2;
		7'd23: data = 3'd0;
		7'd24: data = 3'd5;
		7'd25: data = 3'd3;
		7'd26: data = 3'd1;
		7'd27: data = 3'd0;
		7'd28: data = 3'd5;
		7'd29: data = 3'd3;
		7'd30: data = 3'd2;
		7'd31: data = 3'd0;
		7'd32: data = 3'd3;
		7'd33: data = 3'd3;
		7'd34: data = 3'd1;
		7'd35: data = 3'd0;
		7'd36: data = 3'd6;
		7'd37: data = 3'd3;
		7'd38: data = 3'd1;
		7'd39: data = 3'd0;
		7'd40: data = 3'd6;
		7'd41: data = 3'd4;
		7'd42: data = 3'd1;
		7'd43: data = 3'd0;
		7'd44: data = 3'd2;
		7'd45: data = 3'd2;
		7'd46: data = 3'd0;
		7'd47: data = 3'd0;
		7'd48: data = 3'd6;
		7'd49: data = 3'd3;
		7'd50: data = 3'd2;
		7'd51: data = 3'd0;
		7'd52: data = 3'd2;
		7'd53: data = 3'd0;
		7'd54: data = 3'd0;
		7'd55: data = 3'd0;
		7'd56: data = 3'd0;
		7'd57: data = 3'd0;
		7'd58: data = 3'd1;
		7'd59: data = 3'd1;
		7'd60: data = 3'd1;
		7'd61: data = 3'd0;
		7'd62: data = 3'd1;
		7'd63: data = 3'd1;
		7'd64: data = 3'd1;
		7'd65: data = 3'd0;
		7'd66: data = 3'd1;
		7'd67: data = 3'd0;
		7'd68: data = 3'd0;
		7'd69: data = 3'd0;
		7'd70: data = 3'd0;
		7'd71: data = 3'd1;
		7'd72: data = 3'd0;
		7'd73: data = 3'd1;
		7'd74: data = 3'd1;
		7'd75: data = 3'd0;
		7'd76: data = 3'd4;
		7'd77: data = 3'd4;
		7'd78: data = 3'd2;
		7'd79: data = 3'd0;
		7'd80: data = 3'd1;
		7'd81: data = 3'd2;
		7'd82: data = 3'd1;
		7'd83: data = 3'd0;
		7'd84: data = 3'd2;
		7'd85: data = 3'd2;
		7'd86: data = 3'd2;
		7'd87: data = 3'd0;
		7'd88: data = 3'd2;
		7'd89: data = 3'd1;
		7'd90: data = 3'd0;
		7'd91: data = 3'd1;
		7'd92: data = 3'd1;
		7'd93: data = 3'd0;
		7'd94: data = 3'd0;
		7'd95: data = 3'd1;
		7'd96: data = 3'd0;
		7'd97: data = 3'd0;
		7'd98: data = 3'd1;
		7'd99: data = 3'd0;
		7'd100: data = 3'd3;
		7'd101: data = 3'd2;
		7'd102: data = 3'd2;
		7'd103: data = 3'd0;
		7'd104: data = 3'd0;
		7'd105: data = 3'd1;
		7'd106: data = 3'd1;
		7'd107: data = 3'd1;
		7'd108: data = 3'd7;
		7'd109: data = 3'd4;
		7'd110: data = 3'd2;
		7'd111: data = 3'd0;
		7'd112: data = 3'd7;
		7'd113: data = 3'd5;
		7'd114: data = 3'd2;
		7'd115: data = 3'd0;
		default: data = 3'd0;
	endcase
end
endmodule

module layer1_N0_idx_1(address, data);
input wire [9:0] address;
output reg [4:0] data;

always @(*) begin
	case(address)
		10'd0: data = 5'd0;
		10'd1: data = 5'd0;
		10'd2: data = 5'd5;
		10'd3: data = 5'd14;
		10'd4: data = 5'd0;
		10'd5: data = 5'd0;
		10'd6: data = 5'd1;
		10'd7: data = 5'd15;
		10'd8: data = 5'd0;
		10'd9: data = 5'd5;
		10'd10: data = 5'd1;
		10'd11: data = 5'd15;
		10'd12: data = 5'd0;
		10'd13: data = 5'd0;
		10'd14: data = 5'd0;
		10'd15: data = 5'd16;
		10'd16: data = 5'd0;
		10'd17: data = 5'd3;
		10'd18: data = 5'd0;
		10'd19: data = 5'd0;
		10'd20: data = 5'd0;
		10'd21: data = 5'd0;
		10'd22: data = 5'd2;
		10'd23: data = 5'd0;
		10'd24: data = 5'd0;
		10'd25: data = 5'd0;
		10'd26: data = 5'd1;
		10'd27: data = 5'd3;
		10'd28: data = 5'd5;
		10'd29: data = 5'd0;
		10'd30: data = 5'd1;
		10'd31: data = 5'd8;
		10'd32: data = 5'd3;
		10'd33: data = 5'd1;
		10'd34: data = 5'd0;
		10'd35: data = 5'd0;
		10'd36: data = 5'd5;
		10'd37: data = 5'd0;
		10'd38: data = 5'd1;
		10'd39: data = 5'd2;
		10'd40: data = 5'd3;
		10'd41: data = 5'd2;
		10'd42: data = 5'd3;
		10'd43: data = 5'd2;
		10'd44: data = 5'd3;
		10'd45: data = 5'd1;
		10'd46: data = 5'd2;
		10'd47: data = 5'd4;
		10'd48: data = 5'd5;
		10'd49: data = 5'd3;
		10'd50: data = 5'd0;
		10'd51: data = 5'd4;
		10'd52: data = 5'd0;
		10'd53: data = 5'd2;
		10'd54: data = 5'd0;
		10'd55: data = 5'd1;
		10'd56: data = 5'd0;
		10'd57: data = 5'd0;
		10'd58: data = 5'd5;
		10'd59: data = 5'd1;
		10'd60: data = 5'd0;
		10'd61: data = 5'd1;
		10'd62: data = 5'd0;
		10'd63: data = 5'd7;
		10'd64: data = 5'd0;
		10'd65: data = 5'd0;
		10'd66: data = 5'd2;
		10'd67: data = 5'd14;
		10'd68: data = 5'd0;
		10'd69: data = 5'd5;
		10'd70: data = 5'd3;
		10'd71: data = 5'd17;
		10'd72: data = 5'd0;
		10'd73: data = 5'd3;
		10'd74: data = 5'd3;
		10'd75: data = 5'd0;
		10'd76: data = 5'd0;
		10'd77: data = 5'd3;
		10'd78: data = 5'd0;
		10'd79: data = 5'd5;
		10'd80: data = 5'd0;
		10'd81: data = 5'd1;
		10'd82: data = 5'd2;
		10'd83: data = 5'd0;
		10'd84: data = 5'd0;
		10'd85: data = 5'd0;
		10'd86: data = 5'd1;
		10'd87: data = 5'd11;
		10'd88: data = 5'd0;
		10'd89: data = 5'd0;
		10'd90: data = 5'd0;
		10'd91: data = 5'd0;
		10'd92: data = 5'd21;
		10'd93: data = 5'd0;
		10'd94: data = 5'd0;
		10'd95: data = 5'd0;
		10'd96: data = 5'd3;
		10'd97: data = 5'd0;
		10'd98: data = 5'd0;
		10'd99: data = 5'd8;
		10'd100: data = 5'd5;
		10'd101: data = 5'd3;
		10'd102: data = 5'd0;
		10'd103: data = 5'd1;
		10'd104: data = 5'd11;
		10'd105: data = 5'd2;
		10'd106: data = 5'd2;
		10'd107: data = 5'd2;
		10'd108: data = 5'd3;
		10'd109: data = 5'd1;
		10'd110: data = 5'd0;
		10'd111: data = 5'd2;
		10'd112: data = 5'd5;
		10'd113: data = 5'd3;
		10'd114: data = 5'd0;
		10'd115: data = 5'd7;
		10'd116: data = 5'd0;
		10'd117: data = 5'd2;
		10'd118: data = 5'd0;
		10'd119: data = 5'd1;
		10'd120: data = 5'd0;
		10'd121: data = 5'd1;
		10'd122: data = 5'd1;
		10'd123: data = 5'd1;
		10'd124: data = 5'd0;
		10'd125: data = 5'd3;
		10'd126: data = 5'd0;
		10'd127: data = 5'd7;
		10'd128: data = 5'd0;
		10'd129: data = 5'd5;
		10'd130: data = 5'd22;
		10'd131: data = 5'd0;
		10'd132: data = 5'd0;
		10'd133: data = 5'd3;
		10'd134: data = 5'd1;
		10'd135: data = 5'd0;
		10'd136: data = 5'd0;
		10'd137: data = 5'd2;
		10'd138: data = 5'd3;
		10'd139: data = 5'd18;
		10'd140: data = 5'd0;
		10'd141: data = 5'd0;
		10'd142: data = 5'd0;
		10'd143: data = 5'd5;
		10'd144: data = 5'd0;
		10'd145: data = 5'd0;
		10'd146: data = 5'd2;
		10'd147: data = 5'd1;
		10'd148: data = 5'd0;
		10'd149: data = 5'd2;
		10'd150: data = 5'd1;
		10'd151: data = 5'd0;
		10'd152: data = 5'd5;
		10'd153: data = 5'd0;
		10'd154: data = 5'd9;
		10'd155: data = 5'd4;
		10'd156: data = 5'd3;
		10'd157: data = 5'd2;
		10'd158: data = 5'd0;
		10'd159: data = 5'd0;
		10'd160: data = 5'd5;
		10'd161: data = 5'd3;
		10'd162: data = 5'd0;
		10'd163: data = 5'd2;
		10'd164: data = 5'd8;
		10'd165: data = 5'd3;
		10'd166: data = 5'd2;
		10'd167: data = 5'd2;
		10'd168: data = 5'd11;
		10'd169: data = 5'd2;
		10'd170: data = 5'd0;
		10'd171: data = 5'd0;
		10'd172: data = 5'd3;
		10'd173: data = 5'd0;
		10'd174: data = 5'd2;
		10'd175: data = 5'd1;
		10'd176: data = 5'd5;
		10'd177: data = 5'd3;
		10'd178: data = 5'd0;
		10'd179: data = 5'd2;
		10'd180: data = 5'd0;
		10'd181: data = 5'd1;
		10'd182: data = 5'd0;
		10'd183: data = 5'd3;
		10'd184: data = 5'd0;
		10'd185: data = 5'd0;
		10'd186: data = 5'd0;
		10'd187: data = 5'd1;
		10'd188: data = 5'd0;
		10'd189: data = 5'd2;
		10'd190: data = 5'd0;
		10'd191: data = 5'd7;
		10'd192: data = 5'd0;
		10'd193: data = 5'd3;
		10'd194: data = 5'd0;
		10'd195: data = 5'd14;
		10'd196: data = 5'd0;
		10'd197: data = 5'd1;
		10'd198: data = 5'd1;
		10'd199: data = 5'd0;
		10'd200: data = 5'd0;
		10'd201: data = 5'd0;
		10'd202: data = 5'd0;
		10'd203: data = 5'd5;
		10'd204: data = 5'd0;
		10'd205: data = 5'd8;
		10'd206: data = 5'd2;
		10'd207: data = 5'd0;
		10'd208: data = 5'd0;
		10'd209: data = 5'd0;
		10'd210: data = 5'd0;
		10'd211: data = 5'd1;
		10'd212: data = 5'd0;
		10'd213: data = 5'd0;
		10'd214: data = 5'd1;
		10'd215: data = 5'd0;
		10'd216: data = 5'd5;
		10'd217: data = 5'd0;
		10'd218: data = 5'd1;
		10'd219: data = 5'd2;
		10'd220: data = 5'd3;
		10'd221: data = 5'd0;
		10'd222: data = 5'd0;
		10'd223: data = 5'd0;
		10'd224: data = 5'd8;
		10'd225: data = 5'd3;
		10'd226: data = 5'd0;
		10'd227: data = 5'd8;
		10'd228: data = 5'd8;
		10'd229: data = 5'd1;
		10'd230: data = 5'd0;
		10'd231: data = 5'd19;
		10'd232: data = 5'd11;
		10'd233: data = 5'd0;
		10'd234: data = 5'd2;
		10'd235: data = 5'd2;
		10'd236: data = 5'd3;
		10'd237: data = 5'd3;
		10'd238: data = 5'd0;
		10'd239: data = 5'd0;
		10'd240: data = 5'd5;
		10'd241: data = 5'd0;
		10'd242: data = 5'd2;
		10'd243: data = 5'd1;
		10'd244: data = 5'd5;
		10'd245: data = 5'd0;
		10'd246: data = 5'd0;
		10'd247: data = 5'd2;
		10'd248: data = 5'd0;
		10'd249: data = 5'd2;
		10'd250: data = 5'd0;
		10'd251: data = 5'd3;
		10'd252: data = 5'd0;
		10'd253: data = 5'd0;
		10'd254: data = 5'd0;
		10'd255: data = 5'd2;
		10'd256: data = 5'd0;
		10'd257: data = 5'd0;
		10'd258: data = 5'd23;
		10'd259: data = 5'd0;
		10'd260: data = 5'd0;
		10'd261: data = 5'd1;
		10'd262: data = 5'd0;
		10'd263: data = 5'd5;
		10'd264: data = 5'd0;
		10'd265: data = 5'd0;
		10'd266: data = 5'd2;
		10'd267: data = 5'd20;
		10'd268: data = 5'd0;
		10'd269: data = 5'd0;
		10'd270: data = 5'd0;
		10'd271: data = 5'd0;
		10'd272: data = 5'd5;
		10'd273: data = 5'd5;
		10'd274: data = 5'd5;
		10'd275: data = 5'd2;
		10'd276: data = 5'd5;
		10'd277: data = 5'd0;
		10'd278: data = 5'd2;
		10'd279: data = 5'd0;
		10'd280: data = 5'd0;
		10'd281: data = 5'd0;
		10'd282: data = 5'd0;
		10'd283: data = 5'd0;
		10'd284: data = 5'd3;
		10'd285: data = 5'd0;
		10'd286: data = 5'd0;
		10'd287: data = 5'd0;
		10'd288: data = 5'd8;
		10'd289: data = 5'd0;
		10'd290: data = 5'd0;
		10'd291: data = 5'd1;
		10'd292: data = 5'd0;
		10'd293: data = 5'd0;
		10'd294: data = 5'd2;
		10'd295: data = 5'd1;
		10'd296: data = 5'd0;
		10'd297: data = 5'd2;
		10'd298: data = 5'd0;
		10'd299: data = 5'd19;
		10'd300: data = 5'd2;
		10'd301: data = 5'd0;
		10'd302: data = 5'd2;
		10'd303: data = 5'd2;
		10'd304: data = 5'd3;
		10'd305: data = 5'd0;
		10'd306: data = 5'd0;
		10'd307: data = 5'd0;
		10'd308: data = 5'd5;
		10'd309: data = 5'd2;
		10'd310: data = 5'd0;
		10'd311: data = 5'd1;
		10'd312: data = 5'd0;
		10'd313: data = 5'd0;
		10'd314: data = 5'd0;
		10'd315: data = 5'd3;
		10'd316: data = 5'd0;
		10'd317: data = 5'd3;
		10'd318: data = 5'd0;
		10'd319: data = 5'd1;
		10'd320: data = 5'd0;
		10'd321: data = 5'd1;
		10'd322: data = 5'd0;
		10'd323: data = 5'd24;
		10'd324: data = 5'd0;
		10'd325: data = 5'd0;
		10'd326: data = 5'd1;
		10'd327: data = 5'd5;
		10'd328: data = 5'd5;
		10'd329: data = 5'd9;
		10'd330: data = 5'd0;
		10'd331: data = 5'd0;
		10'd332: data = 5'd5;
		10'd333: data = 5'd0;
		10'd334: data = 5'd0;
		10'd335: data = 5'd1;
		10'd336: data = 5'd5;
		10'd337: data = 5'd0;
		10'd338: data = 5'd2;
		10'd339: data = 5'd2;
		10'd340: data = 5'd3;
		10'd341: data = 5'd0;
		10'd342: data = 5'd12;
		10'd343: data = 5'd0;
		10'd344: data = 5'd3;
		10'd345: data = 5'd0;
		10'd346: data = 5'd0;
		10'd347: data = 5'd0;
		10'd348: data = 5'd3;
		10'd349: data = 5'd0;
		10'd350: data = 5'd4;
		10'd351: data = 5'd0;
		10'd352: data = 5'd8;
		10'd353: data = 5'd0;
		10'd354: data = 5'd0;
		10'd355: data = 5'd10;
		10'd356: data = 5'd0;
		10'd357: data = 5'd0;
		10'd358: data = 5'd0;
		10'd359: data = 5'd10;
		10'd360: data = 5'd0;
		10'd361: data = 5'd0;
		10'd362: data = 5'd2;
		10'd363: data = 5'd1;
		10'd364: data = 5'd0;
		10'd365: data = 5'd0;
		10'd366: data = 5'd0;
		10'd367: data = 5'd8;
		10'd368: data = 5'd3;
		10'd369: data = 5'd0;
		10'd370: data = 5'd3;
		10'd371: data = 5'd1;
		10'd372: data = 5'd0;
		10'd373: data = 5'd0;
		10'd374: data = 5'd0;
		10'd375: data = 5'd8;
		10'd376: data = 5'd5;
		10'd377: data = 5'd3;
		10'd378: data = 5'd0;
		10'd379: data = 5'd2;
		10'd380: data = 5'd0;
		10'd381: data = 5'd0;
		10'd382: data = 5'd0;
		10'd383: data = 5'd1;
		10'd384: data = 5'd5;
		10'd385: data = 5'd2;
		10'd386: data = 5'd17;
		10'd387: data = 5'd5;
		10'd388: data = 5'd5;
		10'd389: data = 5'd0;
		10'd390: data = 5'd1;
		10'd391: data = 5'd3;
		10'd392: data = 5'd5;
		10'd393: data = 5'd0;
		10'd394: data = 5'd0;
		10'd395: data = 5'd0;
		10'd396: data = 5'd0;
		10'd397: data = 5'd2;
		10'd398: data = 5'd2;
		10'd399: data = 5'd1;
		10'd400: data = 5'd3;
		10'd401: data = 5'd0;
		10'd402: data = 5'd0;
		10'd403: data = 5'd2;
		10'd404: data = 5'd3;
		10'd405: data = 5'd0;
		10'd406: data = 5'd1;
		10'd407: data = 5'd0;
		10'd408: data = 5'd11;
		10'd409: data = 5'd0;
		10'd410: data = 5'd4;
		10'd411: data = 5'd2;
		10'd412: data = 5'd8;
		10'd413: data = 5'd0;
		10'd414: data = 5'd4;
		10'd415: data = 5'd2;
		10'd416: data = 5'd8;
		10'd417: data = 5'd0;
		10'd418: data = 5'd1;
		10'd419: data = 5'd1;
		10'd420: data = 5'd0;
		10'd421: data = 5'd0;
		10'd422: data = 5'd2;
		10'd423: data = 5'd1;
		10'd424: data = 5'd0;
		10'd425: data = 5'd0;
		10'd426: data = 5'd0;
		10'd427: data = 5'd10;
		10'd428: data = 5'd0;
		10'd429: data = 5'd0;
		10'd430: data = 5'd2;
		10'd431: data = 5'd1;
		10'd432: data = 5'd1;
		10'd433: data = 5'd0;
		10'd434: data = 5'd0;
		10'd435: data = 5'd8;
		10'd436: data = 5'd3;
		10'd437: data = 5'd0;
		10'd438: data = 5'd3;
		10'd439: data = 5'd2;
		10'd440: data = 5'd5;
		10'd441: data = 5'd0;
		10'd442: data = 5'd0;
		10'd443: data = 5'd1;
		10'd444: data = 5'd5;
		10'd445: data = 5'd0;
		10'd446: data = 5'd0;
		10'd447: data = 5'd2;
		10'd448: data = 5'd5;
		10'd449: data = 5'd0;
		10'd450: data = 5'd0;
		10'd451: data = 5'd5;
		10'd452: data = 5'd5;
		10'd453: data = 5'd9;
		10'd454: data = 5'd0;
		10'd455: data = 5'd3;
		10'd456: data = 5'd3;
		10'd457: data = 5'd0;
		10'd458: data = 5'd1;
		10'd459: data = 5'd1;
		10'd460: data = 5'd3;
		10'd461: data = 5'd0;
		10'd462: data = 5'd0;
		10'd463: data = 5'd2;
		10'd464: data = 5'd3;
		10'd465: data = 5'd0;
		10'd466: data = 5'd2;
		10'd467: data = 5'd2;
		10'd468: data = 5'd0;
		10'd469: data = 5'd0;
		10'd470: data = 5'd1;
		10'd471: data = 5'd9;
		10'd472: data = 5'd0;
		10'd473: data = 5'd0;
		10'd474: data = 5'd4;
		10'd475: data = 5'd0;
		10'd476: data = 5'd0;
		10'd477: data = 5'd2;
		10'd478: data = 5'd1;
		10'd479: data = 5'd0;
		10'd480: data = 5'd0;
		10'd481: data = 5'd1;
		10'd482: data = 5'd1;
		10'd483: data = 5'd1;
		10'd484: data = 5'd0;
		10'd485: data = 5'd4;
		10'd486: data = 5'd2;
		10'd487: data = 5'd1;
		10'd488: data = 5'd0;
		10'd489: data = 5'd1;
		10'd490: data = 5'd25;
		10'd491: data = 5'd1;
		10'd492: data = 5'd0;
		10'd493: data = 5'd0;
		10'd494: data = 5'd0;
		10'd495: data = 5'd0;
		10'd496: data = 5'd0;
		10'd497: data = 5'd0;
		10'd498: data = 5'd3;
		10'd499: data = 5'd2;
		10'd500: data = 5'd2;
		10'd501: data = 5'd0;
		10'd502: data = 5'd0;
		10'd503: data = 5'd8;
		10'd504: data = 5'd3;
		10'd505: data = 5'd0;
		10'd506: data = 5'd0;
		10'd507: data = 5'd2;
		10'd508: data = 5'd5;
		10'd509: data = 5'd0;
		10'd510: data = 5'd1;
		10'd511: data = 5'd1;
		10'd512: data = 5'd3;
		10'd513: data = 5'd1;
		10'd514: data = 5'd0;
		10'd515: data = 5'd3;
		10'd516: data = 5'd3;
		10'd517: data = 5'd0;
		10'd518: data = 5'd1;
		10'd519: data = 5'd0;
		10'd520: data = 5'd3;
		10'd521: data = 5'd0;
		10'd522: data = 5'd0;
		10'd523: data = 5'd1;
		10'd524: data = 5'd0;
		10'd525: data = 5'd0;
		10'd526: data = 5'd2;
		10'd527: data = 5'd2;
		10'd528: data = 5'd0;
		10'd529: data = 5'd0;
		10'd530: data = 5'd2;
		10'd531: data = 5'd13;
		10'd532: data = 5'd0;
		10'd533: data = 5'd0;
		10'd534: data = 5'd12;
		10'd535: data = 5'd0;
		10'd536: data = 5'd1;
		10'd537: data = 5'd0;
		10'd538: data = 5'd1;
		10'd539: data = 5'd1;
		10'd540: data = 5'd2;
		10'd541: data = 5'd2;
		10'd542: data = 5'd1;
		10'd543: data = 5'd1;
		10'd544: data = 5'd0;
		10'd545: data = 5'd7;
		10'd546: data = 5'd2;
		10'd547: data = 5'd0;
		10'd548: data = 5'd0;
		10'd549: data = 5'd0;
		10'd550: data = 5'd0;
		10'd551: data = 5'd0;
		10'd552: data = 5'd0;
		10'd553: data = 5'd0;
		10'd554: data = 5'd2;
		10'd555: data = 5'd1;
		10'd556: data = 5'd12;
		10'd557: data = 5'd0;
		10'd558: data = 5'd2;
		10'd559: data = 5'd1;
		10'd560: data = 5'd0;
		10'd561: data = 5'd0;
		10'd562: data = 5'd0;
		10'd563: data = 5'd0;
		10'd564: data = 5'd0;
		10'd565: data = 5'd0;
		10'd566: data = 5'd3;
		10'd567: data = 5'd2;
		10'd568: data = 5'd3;
		10'd569: data = 5'd0;
		10'd570: data = 5'd0;
		10'd571: data = 5'd1;
		10'd572: data = 5'd0;
		10'd573: data = 5'd0;
		10'd574: data = 5'd0;
		10'd575: data = 5'd2;
		10'd576: data = 5'd3;
		10'd577: data = 5'd12;
		10'd578: data = 5'd0;
		10'd579: data = 5'd3;
		10'd580: data = 5'd0;
		10'd581: data = 5'd1;
		10'd582: data = 5'd15;
		10'd583: data = 5'd0;
		10'd584: data = 5'd0;
		10'd585: data = 5'd0;
		10'd586: data = 5'd1;
		10'd587: data = 5'd2;
		10'd588: data = 5'd0;
		10'd589: data = 5'd0;
		10'd590: data = 5'd2;
		10'd591: data = 5'd2;
		10'd592: data = 5'd1;
		10'd593: data = 5'd0;
		10'd594: data = 5'd3;
		10'd595: data = 5'd1;
		10'd596: data = 5'd1;
		10'd597: data = 5'd0;
		10'd598: data = 5'd0;
		10'd599: data = 5'd1;
		10'd600: data = 5'd1;
		10'd601: data = 5'd2;
		10'd602: data = 5'd10;
		10'd603: data = 5'd1;
		10'd604: data = 5'd1;
		10'd605: data = 5'd4;
		10'd606: data = 5'd10;
		10'd607: data = 5'd0;
		10'd608: data = 5'd2;
		10'd609: data = 5'd1;
		10'd610: data = 5'd0;
		10'd611: data = 5'd0;
		10'd612: data = 5'd0;
		10'd613: data = 5'd2;
		10'd614: data = 5'd4;
		10'd615: data = 5'd0;
		10'd616: data = 5'd2;
		10'd617: data = 5'd0;
		10'd618: data = 5'd0;
		10'd619: data = 5'd0;
		10'd620: data = 5'd4;
		10'd621: data = 5'd0;
		10'd622: data = 5'd0;
		10'd623: data = 5'd1;
		10'd624: data = 5'd4;
		10'd625: data = 5'd0;
		10'd626: data = 5'd3;
		10'd627: data = 5'd9;
		10'd628: data = 5'd0;
		10'd629: data = 5'd0;
		10'd630: data = 5'd0;
		10'd631: data = 5'd1;
		10'd632: data = 5'd0;
		10'd633: data = 5'd0;
		10'd634: data = 5'd0;
		10'd635: data = 5'd2;
		10'd636: data = 5'd3;
		10'd637: data = 5'd0;
		10'd638: data = 5'd1;
		10'd639: data = 5'd2;
		10'd640: data = 5'd0;
		10'd641: data = 5'd0;
		10'd642: data = 5'd0;
		10'd643: data = 5'd0;
		10'd644: data = 5'd0;
		10'd645: data = 5'd0;
		10'd646: data = 5'd0;
		10'd647: data = 5'd1;
		10'd648: data = 5'd4;
		10'd649: data = 5'd0;
		10'd650: data = 5'd2;
		10'd651: data = 5'd2;
		10'd652: data = 5'd4;
		10'd653: data = 5'd0;
		10'd654: data = 5'd3;
		10'd655: data = 5'd1;
		10'd656: data = 5'd4;
		10'd657: data = 5'd0;
		10'd658: data = 5'd0;
		10'd659: data = 5'd2;
		10'd660: data = 5'd7;
		10'd661: data = 5'd0;
		10'd662: data = 5'd0;
		10'd663: data = 5'd1;
		10'd664: data = 5'd6;
		10'd665: data = 5'd2;
		10'd666: data = 5'd10;
		10'd667: data = 5'd0;
		10'd668: data = 5'd7;
		10'd669: data = 5'd4;
		10'd670: data = 5'd0;
		10'd671: data = 5'd0;
		10'd672: data = 5'd1;
		10'd673: data = 5'd1;
		10'd674: data = 5'd0;
		10'd675: data = 5'd0;
		10'd676: data = 5'd2;
		10'd677: data = 5'd7;
		10'd678: data = 5'd1;
		10'd679: data = 5'd0;
		10'd680: data = 5'd1;
		10'd681: data = 5'd1;
		10'd682: data = 5'd4;
		10'd683: data = 5'd0;
		10'd684: data = 5'd4;
		10'd685: data = 5'd0;
		10'd686: data = 5'd0;
		10'd687: data = 5'd0;
		10'd688: data = 5'd4;
		10'd689: data = 5'd0;
		10'd690: data = 5'd0;
		10'd691: data = 5'd13;
		10'd692: data = 5'd4;
		10'd693: data = 5'd0;
		10'd694: data = 5'd0;
		10'd695: data = 5'd10;
		10'd696: data = 5'd0;
		10'd697: data = 5'd0;
		10'd698: data = 5'd0;
		10'd699: data = 5'd1;
		10'd700: data = 5'd2;
		10'd701: data = 5'd0;
		10'd702: data = 5'd0;
		10'd703: data = 5'd0;
		10'd704: data = 5'd4;
		10'd705: data = 5'd1;
		10'd706: data = 5'd26;
		10'd707: data = 5'd0;
		10'd708: data = 5'd4;
		10'd709: data = 5'd0;
		10'd710: data = 5'd16;
		10'd711: data = 5'd1;
		10'd712: data = 5'd4;
		10'd713: data = 5'd0;
		10'd714: data = 5'd0;
		10'd715: data = 5'd2;
		10'd716: data = 5'd6;
		10'd717: data = 5'd0;
		10'd718: data = 5'd0;
		10'd719: data = 5'd0;
		10'd720: data = 5'd6;
		10'd721: data = 5'd0;
		10'd722: data = 5'd0;
		10'd723: data = 5'd1;
		10'd724: data = 5'd6;
		10'd725: data = 5'd2;
		10'd726: data = 5'd0;
		10'd727: data = 5'd0;
		10'd728: data = 5'd6;
		10'd729: data = 5'd4;
		10'd730: data = 5'd0;
		10'd731: data = 5'd0;
		10'd732: data = 5'd6;
		10'd733: data = 5'd4;
		10'd734: data = 5'd1;
		10'd735: data = 5'd0;
		10'd736: data = 5'd6;
		10'd737: data = 5'd6;
		10'd738: data = 5'd9;
		10'd739: data = 5'd0;
		10'd740: data = 5'd1;
		10'd741: data = 5'd1;
		10'd742: data = 5'd10;
		10'd743: data = 5'd0;
		10'd744: data = 5'd1;
		10'd745: data = 5'd7;
		10'd746: data = 5'd4;
		10'd747: data = 5'd0;
		10'd748: data = 5'd4;
		10'd749: data = 5'd4;
		10'd750: data = 5'd0;
		10'd751: data = 5'd0;
		10'd752: data = 5'd4;
		10'd753: data = 5'd1;
		10'd754: data = 5'd0;
		10'd755: data = 5'd1;
		10'd756: data = 5'd4;
		10'd757: data = 5'd0;
		10'd758: data = 5'd0;
		10'd759: data = 5'd1;
		10'd760: data = 5'd4;
		10'd761: data = 5'd0;
		10'd762: data = 5'd0;
		10'd763: data = 5'd10;
		10'd764: data = 5'd0;
		10'd765: data = 5'd0;
		10'd766: data = 5'd1;
		10'd767: data = 5'd1;
		10'd768: data = 5'd4;
		10'd769: data = 5'd0;
		10'd770: data = 5'd0;
		10'd771: data = 5'd1;
		10'd772: data = 5'd1;
		10'd773: data = 5'd1;
		10'd774: data = 5'd5;
		10'd775: data = 5'd2;
		10'd776: data = 5'd4;
		10'd777: data = 5'd0;
		10'd778: data = 5'd1;
		10'd779: data = 5'd1;
		10'd780: data = 5'd4;
		10'd781: data = 5'd0;
		10'd782: data = 5'd0;
		10'd783: data = 5'd0;
		10'd784: data = 5'd7;
		10'd785: data = 5'd0;
		10'd786: data = 5'd0;
		10'd787: data = 5'd0;
		10'd788: data = 5'd6;
		10'd789: data = 5'd0;
		10'd790: data = 5'd0;
		10'd791: data = 5'd0;
		10'd792: data = 5'd6;
		10'd793: data = 5'd4;
		10'd794: data = 5'd1;
		10'd795: data = 5'd0;
		10'd796: data = 5'd6;
		10'd797: data = 5'd1;
		10'd798: data = 5'd1;
		10'd799: data = 5'd0;
		10'd800: data = 5'd0;
		10'd801: data = 5'd7;
		10'd802: data = 5'd1;
		10'd803: data = 5'd0;
		10'd804: data = 5'd7;
		10'd805: data = 5'd1;
		10'd806: data = 5'd1;
		10'd807: data = 5'd0;
		10'd808: data = 5'd1;
		10'd809: data = 5'd1;
		10'd810: data = 5'd10;
		10'd811: data = 5'd0;
		10'd812: data = 5'd4;
		10'd813: data = 5'd2;
		10'd814: data = 5'd4;
		10'd815: data = 5'd0;
		10'd816: data = 5'd4;
		10'd817: data = 5'd0;
		10'd818: data = 5'd0;
		10'd819: data = 5'd0;
		10'd820: data = 5'd4;
		10'd821: data = 5'd0;
		10'd822: data = 5'd4;
		10'd823: data = 5'd1;
		10'd824: data = 5'd4;
		10'd825: data = 5'd0;
		10'd826: data = 5'd0;
		10'd827: data = 5'd1;
		10'd828: data = 5'd1;
		10'd829: data = 5'd1;
		10'd830: data = 5'd0;
		10'd831: data = 5'd0;
		10'd832: data = 5'd4;
		10'd833: data = 5'd1;
		10'd834: data = 5'd18;
		10'd835: data = 5'd1;
		10'd836: data = 5'd4;
		10'd837: data = 5'd0;
		10'd838: data = 5'd2;
		10'd839: data = 5'd1;
		10'd840: data = 5'd6;
		10'd841: data = 5'd0;
		10'd842: data = 5'd1;
		10'd843: data = 5'd0;
		10'd844: data = 5'd6;
		10'd845: data = 5'd0;
		10'd846: data = 5'd0;
		10'd847: data = 5'd0;
		10'd848: data = 5'd6;
		10'd849: data = 5'd0;
		10'd850: data = 5'd0;
		10'd851: data = 5'd0;
		10'd852: data = 5'd6;
		10'd853: data = 5'd4;
		10'd854: data = 5'd1;
		10'd855: data = 5'd0;
		10'd856: data = 5'd0;
		10'd857: data = 5'd4;
		10'd858: data = 5'd1;
		10'd859: data = 5'd0;
		10'd860: data = 5'd0;
		10'd861: data = 5'd1;
		10'd862: data = 5'd1;
		10'd863: data = 5'd0;
		10'd864: data = 5'd0;
		10'd865: data = 5'd7;
		10'd866: data = 5'd1;
		10'd867: data = 5'd0;
		10'd868: data = 5'd0;
		10'd869: data = 5'd7;
		10'd870: data = 5'd13;
		10'd871: data = 5'd0;
		10'd872: data = 5'd6;
		10'd873: data = 5'd1;
		10'd874: data = 5'd1;
		10'd875: data = 5'd0;
		10'd876: data = 5'd7;
		10'd877: data = 5'd7;
		10'd878: data = 5'd10;
		10'd879: data = 5'd0;
		10'd880: data = 5'd7;
		10'd881: data = 5'd1;
		10'd882: data = 5'd4;
		10'd883: data = 5'd0;
		10'd884: data = 5'd6;
		10'd885: data = 5'd0;
		10'd886: data = 5'd4;
		10'd887: data = 5'd0;
		10'd888: data = 5'd6;
		10'd889: data = 5'd1;
		10'd890: data = 5'd1;
		10'd891: data = 5'd1;
		10'd892: data = 5'd4;
		10'd893: data = 5'd0;
		10'd894: data = 5'd0;
		10'd895: data = 5'd1;
		10'd896: data = 5'd6;
		10'd897: data = 5'd2;
		10'd898: data = 5'd5;
		10'd899: data = 5'd2;
		10'd900: data = 5'd1;
		10'd901: data = 5'd0;
		10'd902: data = 5'd0;
		10'd903: data = 5'd1;
		10'd904: data = 5'd4;
		10'd905: data = 5'd0;
		10'd906: data = 5'd1;
		10'd907: data = 5'd0;
		10'd908: data = 5'd7;
		10'd909: data = 5'd0;
		10'd910: data = 5'd0;
		10'd911: data = 5'd0;
		10'd912: data = 5'd9;
		10'd913: data = 5'd0;
		10'd914: data = 5'd1;
		10'd915: data = 5'd0;
		10'd916: data = 5'd6;
		10'd917: data = 5'd4;
		10'd918: data = 5'd1;
		10'd919: data = 5'd0;
		10'd920: data = 5'd6;
		10'd921: data = 5'd1;
		10'd922: data = 5'd0;
		10'd923: data = 5'd0;
		10'd924: data = 5'd27;
		10'd925: data = 5'd6;
		10'd926: data = 5'd0;
		10'd927: data = 5'd0;
		10'd928: data = 5'd9;
		10'd929: data = 5'd1;
		10'd930: data = 5'd0;
		10'd931: data = 5'd0;
		10'd932: data = 5'd0;
		10'd933: data = 5'd7;
		10'd934: data = 5'd1;
		10'd935: data = 5'd0;
		10'd936: data = 5'd0;
		10'd937: data = 5'd7;
		10'd938: data = 5'd13;
		10'd939: data = 5'd0;
		10'd940: data = 5'd6;
		10'd941: data = 5'd1;
		10'd942: data = 5'd1;
		10'd943: data = 5'd0;
		10'd944: data = 5'd6;
		10'd945: data = 5'd7;
		10'd946: data = 5'd9;
		10'd947: data = 5'd0;
		10'd948: data = 5'd4;
		10'd949: data = 5'd1;
		10'd950: data = 5'd4;
		10'd951: data = 5'd0;
		10'd952: data = 5'd4;
		10'd953: data = 5'd0;
		10'd954: data = 5'd1;
		10'd955: data = 5'd0;
		10'd956: data = 5'd4;
		10'd957: data = 5'd1;
		10'd958: data = 5'd1;
		10'd959: data = 5'd1;
		10'd960: data = 5'd4;
		10'd961: data = 5'd0;
		10'd962: data = 5'd20;
		10'd963: data = 5'd1;
		10'd964: data = 5'd6;
		10'd965: data = 5'd1;
		10'd966: data = 5'd0;
		10'd967: data = 5'd0;
		10'd968: data = 5'd6;
		10'd969: data = 5'd0;
		10'd970: data = 5'd9;
		10'd971: data = 5'd1;
		10'd972: data = 5'd6;
		10'd973: data = 5'd0;
		10'd974: data = 5'd11;
		10'd975: data = 5'd0;
		10'd976: data = 5'd6;
		10'd977: data = 5'd4;
		10'd978: data = 5'd1;
		10'd979: data = 5'd0;
		10'd980: data = 5'd0;
		10'd981: data = 5'd1;
		10'd982: data = 5'd1;
		10'd983: data = 5'd0;
		10'd984: data = 5'd0;
		10'd985: data = 5'd1;
		10'd986: data = 5'd0;
		10'd987: data = 5'd0;
		10'd988: data = 5'd28;
		10'd989: data = 5'd7;
		10'd990: data = 5'd0;
		10'd991: data = 5'd0;
		10'd992: data = 5'd10;
		10'd993: data = 5'd1;
		10'd994: data = 5'd0;
		10'd995: data = 5'd0;
		10'd996: data = 5'd9;
		10'd997: data = 5'd1;
		10'd998: data = 5'd0;
		10'd999: data = 5'd0;
		10'd1000: data = 5'd0;
		10'd1001: data = 5'd7;
		10'd1002: data = 5'd1;
		10'd1003: data = 5'd0;
		10'd1004: data = 5'd12;
		10'd1005: data = 5'd6;
		10'd1006: data = 5'd1;
		10'd1007: data = 5'd0;
		10'd1008: data = 5'd0;
		10'd1009: data = 5'd7;
		10'd1010: data = 5'd1;
		10'd1011: data = 5'd0;
		10'd1012: data = 5'd4;
		10'd1013: data = 5'd2;
		10'd1014: data = 5'd9;
		10'd1015: data = 5'd0;
		10'd1016: data = 5'd4;
		10'd1017: data = 5'd1;
		10'd1018: data = 5'd1;
		10'd1019: data = 5'd0;
		10'd1020: data = 5'd4;
		10'd1021: data = 5'd0;
		10'd1022: data = 5'd2;
		10'd1023: data = 5'd0;
		default: data = 5'd0;
	endcase
end
endmodule

module layer1_N0_rsh_1(address, data);
input wire [9:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		10'd0: data = 2'd3;
		10'd1: data = 2'd3;
		10'd2: data = 2'd1;
		10'd3: data = 2'd0;
		10'd4: data = 2'd3;
		10'd5: data = 2'd3;
		10'd6: data = 2'd2;
		10'd7: data = 2'd0;
		10'd8: data = 2'd3;
		10'd9: data = 2'd1;
		10'd10: data = 2'd2;
		10'd11: data = 2'd0;
		10'd12: data = 2'd3;
		10'd13: data = 2'd2;
		10'd14: data = 2'd2;
		10'd15: data = 2'd0;
		10'd16: data = 2'd3;
		10'd17: data = 2'd1;
		10'd18: data = 2'd2;
		10'd19: data = 2'd1;
		10'd20: data = 2'd3;
		10'd21: data = 2'd1;
		10'd22: data = 2'd1;
		10'd23: data = 2'd1;
		10'd24: data = 2'd3;
		10'd25: data = 2'd1;
		10'd26: data = 2'd1;
		10'd27: data = 2'd1;
		10'd28: data = 2'd1;
		10'd29: data = 2'd1;
		10'd30: data = 2'd1;
		10'd31: data = 2'd0;
		10'd32: data = 2'd1;
		10'd33: data = 2'd1;
		10'd34: data = 2'd1;
		10'd35: data = 2'd1;
		10'd36: data = 2'd0;
		10'd37: data = 2'd1;
		10'd38: data = 2'd1;
		10'd39: data = 2'd0;
		10'd40: data = 2'd1;
		10'd41: data = 2'd1;
		10'd42: data = 2'd1;
		10'd43: data = 2'd0;
		10'd44: data = 2'd1;
		10'd45: data = 2'd1;
		10'd46: data = 2'd1;
		10'd47: data = 2'd0;
		10'd48: data = 2'd1;
		10'd49: data = 2'd1;
		10'd50: data = 2'd1;
		10'd51: data = 2'd0;
		10'd52: data = 2'd3;
		10'd53: data = 2'd1;
		10'd54: data = 2'd1;
		10'd55: data = 2'd0;
		10'd56: data = 2'd3;
		10'd57: data = 2'd1;
		10'd58: data = 2'd0;
		10'd59: data = 2'd0;
		10'd60: data = 2'd3;
		10'd61: data = 2'd1;
		10'd62: data = 2'd1;
		10'd63: data = 2'd0;
		10'd64: data = 2'd3;
		10'd65: data = 2'd3;
		10'd66: data = 2'd1;
		10'd67: data = 2'd0;
		10'd68: data = 2'd3;
		10'd69: data = 2'd1;
		10'd70: data = 2'd1;
		10'd71: data = 2'd0;
		10'd72: data = 2'd3;
		10'd73: data = 2'd1;
		10'd74: data = 2'd1;
		10'd75: data = 2'd3;
		10'd76: data = 2'd3;
		10'd77: data = 2'd1;
		10'd78: data = 2'd2;
		10'd79: data = 2'd1;
		10'd80: data = 2'd3;
		10'd81: data = 2'd1;
		10'd82: data = 2'd1;
		10'd83: data = 2'd2;
		10'd84: data = 2'd3;
		10'd85: data = 2'd1;
		10'd86: data = 2'd1;
		10'd87: data = 2'd0;
		10'd88: data = 2'd3;
		10'd89: data = 2'd1;
		10'd90: data = 2'd1;
		10'd91: data = 2'd1;
		10'd92: data = 2'd0;
		10'd93: data = 2'd1;
		10'd94: data = 2'd1;
		10'd95: data = 2'd1;
		10'd96: data = 2'd1;
		10'd97: data = 2'd1;
		10'd98: data = 2'd1;
		10'd99: data = 2'd0;
		10'd100: data = 2'd0;
		10'd101: data = 2'd1;
		10'd102: data = 2'd1;
		10'd103: data = 2'd0;
		10'd104: data = 2'd0;
		10'd105: data = 2'd1;
		10'd106: data = 2'd1;
		10'd107: data = 2'd0;
		10'd108: data = 2'd1;
		10'd109: data = 2'd1;
		10'd110: data = 2'd1;
		10'd111: data = 2'd0;
		10'd112: data = 2'd1;
		10'd113: data = 2'd1;
		10'd114: data = 2'd1;
		10'd115: data = 2'd0;
		10'd116: data = 2'd3;
		10'd117: data = 2'd1;
		10'd118: data = 2'd1;
		10'd119: data = 2'd0;
		10'd120: data = 2'd3;
		10'd121: data = 2'd1;
		10'd122: data = 2'd0;
		10'd123: data = 2'd0;
		10'd124: data = 2'd3;
		10'd125: data = 2'd1;
		10'd126: data = 2'd1;
		10'd127: data = 2'd0;
		10'd128: data = 2'd3;
		10'd129: data = 2'd1;
		10'd130: data = 2'd0;
		10'd131: data = 2'd3;
		10'd132: data = 2'd3;
		10'd133: data = 2'd1;
		10'd134: data = 2'd1;
		10'd135: data = 2'd3;
		10'd136: data = 2'd3;
		10'd137: data = 2'd1;
		10'd138: data = 2'd1;
		10'd139: data = 2'd0;
		10'd140: data = 2'd3;
		10'd141: data = 2'd1;
		10'd142: data = 2'd2;
		10'd143: data = 2'd1;
		10'd144: data = 2'd3;
		10'd145: data = 2'd1;
		10'd146: data = 2'd1;
		10'd147: data = 2'd1;
		10'd148: data = 2'd3;
		10'd149: data = 2'd1;
		10'd150: data = 2'd2;
		10'd151: data = 2'd1;
		10'd152: data = 2'd1;
		10'd153: data = 2'd1;
		10'd154: data = 2'd1;
		10'd155: data = 2'd0;
		10'd156: data = 2'd1;
		10'd157: data = 2'd1;
		10'd158: data = 2'd1;
		10'd159: data = 2'd1;
		10'd160: data = 2'd0;
		10'd161: data = 2'd1;
		10'd162: data = 2'd1;
		10'd163: data = 2'd0;
		10'd164: data = 2'd0;
		10'd165: data = 2'd1;
		10'd166: data = 2'd1;
		10'd167: data = 2'd0;
		10'd168: data = 2'd0;
		10'd169: data = 2'd1;
		10'd170: data = 2'd1;
		10'd171: data = 2'd1;
		10'd172: data = 2'd1;
		10'd173: data = 2'd1;
		10'd174: data = 2'd1;
		10'd175: data = 2'd0;
		10'd176: data = 2'd1;
		10'd177: data = 2'd1;
		10'd178: data = 2'd1;
		10'd179: data = 2'd0;
		10'd180: data = 2'd3;
		10'd181: data = 2'd1;
		10'd182: data = 2'd1;
		10'd183: data = 2'd0;
		10'd184: data = 2'd3;
		10'd185: data = 2'd1;
		10'd186: data = 2'd1;
		10'd187: data = 2'd0;
		10'd188: data = 2'd3;
		10'd189: data = 2'd1;
		10'd190: data = 2'd1;
		10'd191: data = 2'd0;
		10'd192: data = 2'd3;
		10'd193: data = 2'd1;
		10'd194: data = 2'd3;
		10'd195: data = 2'd0;
		10'd196: data = 2'd3;
		10'd197: data = 2'd1;
		10'd198: data = 2'd2;
		10'd199: data = 2'd3;
		10'd200: data = 2'd3;
		10'd201: data = 2'd1;
		10'd202: data = 2'd2;
		10'd203: data = 2'd1;
		10'd204: data = 2'd3;
		10'd205: data = 2'd0;
		10'd206: data = 2'd1;
		10'd207: data = 2'd2;
		10'd208: data = 2'd3;
		10'd209: data = 2'd1;
		10'd210: data = 2'd2;
		10'd211: data = 2'd1;
		10'd212: data = 2'd3;
		10'd213: data = 2'd1;
		10'd214: data = 2'd1;
		10'd215: data = 2'd1;
		10'd216: data = 2'd1;
		10'd217: data = 2'd1;
		10'd218: data = 2'd1;
		10'd219: data = 2'd0;
		10'd220: data = 2'd1;
		10'd221: data = 2'd1;
		10'd222: data = 2'd1;
		10'd223: data = 2'd1;
		10'd224: data = 2'd0;
		10'd225: data = 2'd1;
		10'd226: data = 2'd1;
		10'd227: data = 2'd0;
		10'd228: data = 2'd0;
		10'd229: data = 2'd1;
		10'd230: data = 2'd1;
		10'd231: data = 2'd0;
		10'd232: data = 2'd0;
		10'd233: data = 2'd1;
		10'd234: data = 2'd1;
		10'd235: data = 2'd0;
		10'd236: data = 2'd1;
		10'd237: data = 2'd1;
		10'd238: data = 2'd1;
		10'd239: data = 2'd1;
		10'd240: data = 2'd1;
		10'd241: data = 2'd1;
		10'd242: data = 2'd1;
		10'd243: data = 2'd0;
		10'd244: data = 2'd1;
		10'd245: data = 2'd1;
		10'd246: data = 2'd1;
		10'd247: data = 2'd0;
		10'd248: data = 2'd3;
		10'd249: data = 2'd1;
		10'd250: data = 2'd1;
		10'd251: data = 2'd0;
		10'd252: data = 2'd3;
		10'd253: data = 2'd1;
		10'd254: data = 2'd1;
		10'd255: data = 2'd0;
		10'd256: data = 2'd3;
		10'd257: data = 2'd1;
		10'd258: data = 2'd0;
		10'd259: data = 2'd3;
		10'd260: data = 2'd3;
		10'd261: data = 2'd1;
		10'd262: data = 2'd2;
		10'd263: data = 2'd1;
		10'd264: data = 2'd3;
		10'd265: data = 2'd1;
		10'd266: data = 2'd1;
		10'd267: data = 2'd0;
		10'd268: data = 2'd3;
		10'd269: data = 2'd1;
		10'd270: data = 2'd2;
		10'd271: data = 2'd2;
		10'd272: data = 2'd1;
		10'd273: data = 2'd0;
		10'd274: data = 2'd1;
		10'd275: data = 2'd1;
		10'd276: data = 2'd1;
		10'd277: data = 2'd1;
		10'd278: data = 2'd1;
		10'd279: data = 2'd1;
		10'd280: data = 2'd2;
		10'd281: data = 2'd1;
		10'd282: data = 2'd1;
		10'd283: data = 2'd1;
		10'd284: data = 2'd1;
		10'd285: data = 2'd1;
		10'd286: data = 2'd1;
		10'd287: data = 2'd1;
		10'd288: data = 2'd0;
		10'd289: data = 2'd1;
		10'd290: data = 2'd1;
		10'd291: data = 2'd0;
		10'd292: data = 2'd1;
		10'd293: data = 2'd1;
		10'd294: data = 2'd1;
		10'd295: data = 2'd0;
		10'd296: data = 2'd1;
		10'd297: data = 2'd1;
		10'd298: data = 2'd1;
		10'd299: data = 2'd0;
		10'd300: data = 2'd1;
		10'd301: data = 2'd1;
		10'd302: data = 2'd1;
		10'd303: data = 2'd0;
		10'd304: data = 2'd1;
		10'd305: data = 2'd1;
		10'd306: data = 2'd1;
		10'd307: data = 2'd1;
		10'd308: data = 2'd1;
		10'd309: data = 2'd1;
		10'd310: data = 2'd1;
		10'd311: data = 2'd0;
		10'd312: data = 2'd3;
		10'd313: data = 2'd1;
		10'd314: data = 2'd1;
		10'd315: data = 2'd0;
		10'd316: data = 2'd3;
		10'd317: data = 2'd1;
		10'd318: data = 2'd1;
		10'd319: data = 2'd0;
		10'd320: data = 2'd3;
		10'd321: data = 2'd1;
		10'd322: data = 2'd3;
		10'd323: data = 2'd0;
		10'd324: data = 2'd3;
		10'd325: data = 2'd1;
		10'd326: data = 2'd2;
		10'd327: data = 2'd1;
		10'd328: data = 2'd1;
		10'd329: data = 2'd1;
		10'd330: data = 2'd2;
		10'd331: data = 2'd2;
		10'd332: data = 2'd1;
		10'd333: data = 2'd1;
		10'd334: data = 2'd2;
		10'd335: data = 2'd1;
		10'd336: data = 2'd1;
		10'd337: data = 2'd1;
		10'd338: data = 2'd1;
		10'd339: data = 2'd1;
		10'd340: data = 2'd1;
		10'd341: data = 2'd1;
		10'd342: data = 2'd1;
		10'd343: data = 2'd1;
		10'd344: data = 2'd1;
		10'd345: data = 2'd1;
		10'd346: data = 2'd1;
		10'd347: data = 2'd1;
		10'd348: data = 2'd1;
		10'd349: data = 2'd1;
		10'd350: data = 2'd0;
		10'd351: data = 2'd1;
		10'd352: data = 2'd0;
		10'd353: data = 2'd1;
		10'd354: data = 2'd1;
		10'd355: data = 2'd1;
		10'd356: data = 2'd1;
		10'd357: data = 2'd1;
		10'd358: data = 2'd1;
		10'd359: data = 2'd1;
		10'd360: data = 2'd1;
		10'd361: data = 2'd1;
		10'd362: data = 2'd1;
		10'd363: data = 2'd0;
		10'd364: data = 2'd1;
		10'd365: data = 2'd1;
		10'd366: data = 2'd1;
		10'd367: data = 2'd0;
		10'd368: data = 2'd1;
		10'd369: data = 2'd1;
		10'd370: data = 2'd1;
		10'd371: data = 2'd0;
		10'd372: data = 2'd2;
		10'd373: data = 2'd1;
		10'd374: data = 2'd1;
		10'd375: data = 2'd0;
		10'd376: data = 2'd1;
		10'd377: data = 2'd1;
		10'd378: data = 2'd1;
		10'd379: data = 2'd0;
		10'd380: data = 2'd3;
		10'd381: data = 2'd1;
		10'd382: data = 2'd1;
		10'd383: data = 2'd0;
		10'd384: data = 2'd1;
		10'd385: data = 2'd1;
		10'd386: data = 2'd0;
		10'd387: data = 2'd1;
		10'd388: data = 2'd1;
		10'd389: data = 2'd1;
		10'd390: data = 2'd2;
		10'd391: data = 2'd1;
		10'd392: data = 2'd1;
		10'd393: data = 2'd1;
		10'd394: data = 2'd2;
		10'd395: data = 2'd2;
		10'd396: data = 2'd2;
		10'd397: data = 2'd0;
		10'd398: data = 2'd1;
		10'd399: data = 2'd1;
		10'd400: data = 2'd1;
		10'd401: data = 2'd1;
		10'd402: data = 2'd2;
		10'd403: data = 2'd1;
		10'd404: data = 2'd1;
		10'd405: data = 2'd1;
		10'd406: data = 2'd1;
		10'd407: data = 2'd1;
		10'd408: data = 2'd0;
		10'd409: data = 2'd1;
		10'd410: data = 2'd0;
		10'd411: data = 2'd1;
		10'd412: data = 2'd0;
		10'd413: data = 2'd1;
		10'd414: data = 2'd0;
		10'd415: data = 2'd1;
		10'd416: data = 2'd0;
		10'd417: data = 2'd1;
		10'd418: data = 2'd0;
		10'd419: data = 2'd1;
		10'd420: data = 2'd1;
		10'd421: data = 2'd1;
		10'd422: data = 2'd0;
		10'd423: data = 2'd1;
		10'd424: data = 2'd1;
		10'd425: data = 2'd1;
		10'd426: data = 2'd1;
		10'd427: data = 2'd1;
		10'd428: data = 2'd1;
		10'd429: data = 2'd1;
		10'd430: data = 2'd1;
		10'd431: data = 2'd0;
		10'd432: data = 2'd1;
		10'd433: data = 2'd1;
		10'd434: data = 2'd1;
		10'd435: data = 2'd0;
		10'd436: data = 2'd1;
		10'd437: data = 2'd1;
		10'd438: data = 2'd1;
		10'd439: data = 2'd0;
		10'd440: data = 2'd1;
		10'd441: data = 2'd1;
		10'd442: data = 2'd1;
		10'd443: data = 2'd0;
		10'd444: data = 2'd1;
		10'd445: data = 2'd1;
		10'd446: data = 2'd1;
		10'd447: data = 2'd0;
		10'd448: data = 2'd1;
		10'd449: data = 2'd1;
		10'd450: data = 2'd3;
		10'd451: data = 2'd1;
		10'd452: data = 2'd1;
		10'd453: data = 2'd1;
		10'd454: data = 2'd3;
		10'd455: data = 2'd1;
		10'd456: data = 2'd1;
		10'd457: data = 2'd1;
		10'd458: data = 2'd2;
		10'd459: data = 2'd1;
		10'd460: data = 2'd1;
		10'd461: data = 2'd1;
		10'd462: data = 2'd2;
		10'd463: data = 2'd1;
		10'd464: data = 2'd1;
		10'd465: data = 2'd1;
		10'd466: data = 2'd1;
		10'd467: data = 2'd1;
		10'd468: data = 2'd1;
		10'd469: data = 2'd1;
		10'd470: data = 2'd1;
		10'd471: data = 2'd1;
		10'd472: data = 2'd1;
		10'd473: data = 2'd1;
		10'd474: data = 2'd0;
		10'd475: data = 2'd1;
		10'd476: data = 2'd1;
		10'd477: data = 2'd0;
		10'd478: data = 2'd0;
		10'd479: data = 2'd2;
		10'd480: data = 2'd1;
		10'd481: data = 2'd0;
		10'd482: data = 2'd0;
		10'd483: data = 2'd2;
		10'd484: data = 2'd1;
		10'd485: data = 2'd0;
		10'd486: data = 2'd0;
		10'd487: data = 2'd2;
		10'd488: data = 2'd1;
		10'd489: data = 2'd0;
		10'd490: data = 2'd0;
		10'd491: data = 2'd1;
		10'd492: data = 2'd1;
		10'd493: data = 2'd1;
		10'd494: data = 2'd1;
		10'd495: data = 2'd1;
		10'd496: data = 2'd1;
		10'd497: data = 2'd1;
		10'd498: data = 2'd1;
		10'd499: data = 2'd0;
		10'd500: data = 2'd1;
		10'd501: data = 2'd1;
		10'd502: data = 2'd1;
		10'd503: data = 2'd0;
		10'd504: data = 2'd1;
		10'd505: data = 2'd1;
		10'd506: data = 2'd1;
		10'd507: data = 2'd0;
		10'd508: data = 2'd1;
		10'd509: data = 2'd1;
		10'd510: data = 2'd1;
		10'd511: data = 2'd0;
		10'd512: data = 2'd1;
		10'd513: data = 2'd1;
		10'd514: data = 2'd3;
		10'd515: data = 2'd1;
		10'd516: data = 2'd1;
		10'd517: data = 2'd1;
		10'd518: data = 2'd2;
		10'd519: data = 2'd2;
		10'd520: data = 2'd1;
		10'd521: data = 2'd1;
		10'd522: data = 2'd2;
		10'd523: data = 2'd1;
		10'd524: data = 2'd1;
		10'd525: data = 2'd1;
		10'd526: data = 2'd1;
		10'd527: data = 2'd1;
		10'd528: data = 2'd1;
		10'd529: data = 2'd1;
		10'd530: data = 2'd1;
		10'd531: data = 2'd0;
		10'd532: data = 2'd1;
		10'd533: data = 2'd1;
		10'd534: data = 2'd1;
		10'd535: data = 2'd1;
		10'd536: data = 2'd0;
		10'd537: data = 2'd1;
		10'd538: data = 2'd0;
		10'd539: data = 2'd1;
		10'd540: data = 2'd0;
		10'd541: data = 2'd0;
		10'd542: data = 2'd0;
		10'd543: data = 2'd2;
		10'd544: data = 2'd1;
		10'd545: data = 2'd0;
		10'd546: data = 2'd0;
		10'd547: data = 2'd3;
		10'd548: data = 2'd1;
		10'd549: data = 2'd1;
		10'd550: data = 2'd1;
		10'd551: data = 2'd3;
		10'd552: data = 2'd1;
		10'd553: data = 2'd1;
		10'd554: data = 2'd0;
		10'd555: data = 2'd2;
		10'd556: data = 2'd1;
		10'd557: data = 2'd1;
		10'd558: data = 2'd1;
		10'd559: data = 2'd1;
		10'd560: data = 2'd1;
		10'd561: data = 2'd1;
		10'd562: data = 2'd1;
		10'd563: data = 2'd1;
		10'd564: data = 2'd1;
		10'd565: data = 2'd1;
		10'd566: data = 2'd1;
		10'd567: data = 2'd0;
		10'd568: data = 2'd1;
		10'd569: data = 2'd1;
		10'd570: data = 2'd1;
		10'd571: data = 2'd0;
		10'd572: data = 2'd2;
		10'd573: data = 2'd1;
		10'd574: data = 2'd1;
		10'd575: data = 2'd0;
		10'd576: data = 2'd1;
		10'd577: data = 2'd1;
		10'd578: data = 2'd3;
		10'd579: data = 2'd1;
		10'd580: data = 2'd1;
		10'd581: data = 2'd1;
		10'd582: data = 2'd0;
		10'd583: data = 2'd2;
		10'd584: data = 2'd1;
		10'd585: data = 2'd1;
		10'd586: data = 2'd1;
		10'd587: data = 2'd1;
		10'd588: data = 2'd1;
		10'd589: data = 2'd1;
		10'd590: data = 2'd1;
		10'd591: data = 2'd1;
		10'd592: data = 2'd0;
		10'd593: data = 2'd1;
		10'd594: data = 2'd1;
		10'd595: data = 2'd1;
		10'd596: data = 2'd0;
		10'd597: data = 2'd1;
		10'd598: data = 2'd1;
		10'd599: data = 2'd1;
		10'd600: data = 2'd0;
		10'd601: data = 2'd0;
		10'd602: data = 2'd1;
		10'd603: data = 2'd2;
		10'd604: data = 2'd0;
		10'd605: data = 2'd0;
		10'd606: data = 2'd1;
		10'd607: data = 2'd3;
		10'd608: data = 2'd0;
		10'd609: data = 2'd0;
		10'd610: data = 2'd1;
		10'd611: data = 2'd3;
		10'd612: data = 2'd1;
		10'd613: data = 2'd0;
		10'd614: data = 2'd0;
		10'd615: data = 2'd3;
		10'd616: data = 2'd0;
		10'd617: data = 2'd1;
		10'd618: data = 2'd1;
		10'd619: data = 2'd3;
		10'd620: data = 2'd0;
		10'd621: data = 2'd1;
		10'd622: data = 2'd1;
		10'd623: data = 2'd2;
		10'd624: data = 2'd0;
		10'd625: data = 2'd1;
		10'd626: data = 2'd1;
		10'd627: data = 2'd1;
		10'd628: data = 2'd1;
		10'd629: data = 2'd1;
		10'd630: data = 2'd1;
		10'd631: data = 2'd0;
		10'd632: data = 2'd1;
		10'd633: data = 2'd1;
		10'd634: data = 2'd1;
		10'd635: data = 2'd0;
		10'd636: data = 2'd1;
		10'd637: data = 2'd1;
		10'd638: data = 2'd1;
		10'd639: data = 2'd0;
		10'd640: data = 2'd1;
		10'd641: data = 2'd1;
		10'd642: data = 2'd3;
		10'd643: data = 2'd2;
		10'd644: data = 2'd1;
		10'd645: data = 2'd1;
		10'd646: data = 2'd3;
		10'd647: data = 2'd1;
		10'd648: data = 2'd0;
		10'd649: data = 2'd1;
		10'd650: data = 2'd1;
		10'd651: data = 2'd1;
		10'd652: data = 2'd0;
		10'd653: data = 2'd1;
		10'd654: data = 2'd1;
		10'd655: data = 2'd2;
		10'd656: data = 2'd0;
		10'd657: data = 2'd1;
		10'd658: data = 2'd1;
		10'd659: data = 2'd1;
		10'd660: data = 2'd0;
		10'd661: data = 2'd1;
		10'd662: data = 2'd1;
		10'd663: data = 2'd2;
		10'd664: data = 2'd0;
		10'd665: data = 2'd0;
		10'd666: data = 2'd1;
		10'd667: data = 2'd3;
		10'd668: data = 2'd0;
		10'd669: data = 2'd0;
		10'd670: data = 2'd1;
		10'd671: data = 2'd3;
		10'd672: data = 2'd0;
		10'd673: data = 2'd0;
		10'd674: data = 2'd1;
		10'd675: data = 2'd3;
		10'd676: data = 2'd0;
		10'd677: data = 2'd0;
		10'd678: data = 2'd0;
		10'd679: data = 2'd3;
		10'd680: data = 2'd0;
		10'd681: data = 2'd0;
		10'd682: data = 2'd0;
		10'd683: data = 2'd3;
		10'd684: data = 2'd0;
		10'd685: data = 2'd1;
		10'd686: data = 2'd1;
		10'd687: data = 2'd3;
		10'd688: data = 2'd0;
		10'd689: data = 2'd1;
		10'd690: data = 2'd1;
		10'd691: data = 2'd0;
		10'd692: data = 2'd0;
		10'd693: data = 2'd1;
		10'd694: data = 2'd1;
		10'd695: data = 2'd1;
		10'd696: data = 2'd1;
		10'd697: data = 2'd1;
		10'd698: data = 2'd1;
		10'd699: data = 2'd0;
		10'd700: data = 2'd1;
		10'd701: data = 2'd1;
		10'd702: data = 2'd1;
		10'd703: data = 2'd1;
		10'd704: data = 2'd0;
		10'd705: data = 2'd1;
		10'd706: data = 2'd0;
		10'd707: data = 2'd2;
		10'd708: data = 2'd0;
		10'd709: data = 2'd1;
		10'd710: data = 2'd0;
		10'd711: data = 2'd1;
		10'd712: data = 2'd0;
		10'd713: data = 2'd1;
		10'd714: data = 2'd2;
		10'd715: data = 2'd1;
		10'd716: data = 2'd0;
		10'd717: data = 2'd1;
		10'd718: data = 2'd1;
		10'd719: data = 2'd2;
		10'd720: data = 2'd0;
		10'd721: data = 2'd1;
		10'd722: data = 2'd1;
		10'd723: data = 2'd2;
		10'd724: data = 2'd0;
		10'd725: data = 2'd0;
		10'd726: data = 2'd1;
		10'd727: data = 2'd3;
		10'd728: data = 2'd0;
		10'd729: data = 2'd0;
		10'd730: data = 2'd1;
		10'd731: data = 2'd3;
		10'd732: data = 2'd0;
		10'd733: data = 2'd0;
		10'd734: data = 2'd1;
		10'd735: data = 2'd3;
		10'd736: data = 2'd0;
		10'd737: data = 2'd0;
		10'd738: data = 2'd1;
		10'd739: data = 2'd3;
		10'd740: data = 2'd0;
		10'd741: data = 2'd0;
		10'd742: data = 2'd1;
		10'd743: data = 2'd3;
		10'd744: data = 2'd0;
		10'd745: data = 2'd0;
		10'd746: data = 2'd0;
		10'd747: data = 2'd3;
		10'd748: data = 2'd0;
		10'd749: data = 2'd0;
		10'd750: data = 2'd1;
		10'd751: data = 2'd3;
		10'd752: data = 2'd0;
		10'd753: data = 2'd0;
		10'd754: data = 2'd1;
		10'd755: data = 2'd2;
		10'd756: data = 2'd0;
		10'd757: data = 2'd1;
		10'd758: data = 2'd1;
		10'd759: data = 2'd1;
		10'd760: data = 2'd0;
		10'd761: data = 2'd1;
		10'd762: data = 2'd1;
		10'd763: data = 2'd1;
		10'd764: data = 2'd1;
		10'd765: data = 2'd1;
		10'd766: data = 2'd1;
		10'd767: data = 2'd0;
		10'd768: data = 2'd0;
		10'd769: data = 2'd1;
		10'd770: data = 2'd3;
		10'd771: data = 2'd1;
		10'd772: data = 2'd0;
		10'd773: data = 2'd1;
		10'd774: data = 2'd1;
		10'd775: data = 2'd1;
		10'd776: data = 2'd0;
		10'd777: data = 2'd1;
		10'd778: data = 2'd1;
		10'd779: data = 2'd2;
		10'd780: data = 2'd0;
		10'd781: data = 2'd1;
		10'd782: data = 2'd1;
		10'd783: data = 2'd3;
		10'd784: data = 2'd0;
		10'd785: data = 2'd1;
		10'd786: data = 2'd1;
		10'd787: data = 2'd3;
		10'd788: data = 2'd0;
		10'd789: data = 2'd1;
		10'd790: data = 2'd1;
		10'd791: data = 2'd3;
		10'd792: data = 2'd0;
		10'd793: data = 2'd0;
		10'd794: data = 2'd1;
		10'd795: data = 2'd3;
		10'd796: data = 2'd0;
		10'd797: data = 2'd0;
		10'd798: data = 2'd2;
		10'd799: data = 2'd3;
		10'd800: data = 2'd0;
		10'd801: data = 2'd0;
		10'd802: data = 2'd1;
		10'd803: data = 2'd3;
		10'd804: data = 2'd0;
		10'd805: data = 2'd0;
		10'd806: data = 2'd1;
		10'd807: data = 2'd3;
		10'd808: data = 2'd0;
		10'd809: data = 2'd0;
		10'd810: data = 2'd1;
		10'd811: data = 2'd3;
		10'd812: data = 2'd0;
		10'd813: data = 2'd0;
		10'd814: data = 2'd0;
		10'd815: data = 2'd3;
		10'd816: data = 2'd0;
		10'd817: data = 2'd1;
		10'd818: data = 2'd1;
		10'd819: data = 2'd3;
		10'd820: data = 2'd0;
		10'd821: data = 2'd1;
		10'd822: data = 2'd0;
		10'd823: data = 2'd2;
		10'd824: data = 2'd0;
		10'd825: data = 2'd1;
		10'd826: data = 2'd1;
		10'd827: data = 2'd1;
		10'd828: data = 2'd0;
		10'd829: data = 2'd1;
		10'd830: data = 2'd1;
		10'd831: data = 2'd1;
		10'd832: data = 2'd0;
		10'd833: data = 2'd1;
		10'd834: data = 2'd0;
		10'd835: data = 2'd1;
		10'd836: data = 2'd0;
		10'd837: data = 2'd1;
		10'd838: data = 2'd1;
		10'd839: data = 2'd2;
		10'd840: data = 2'd0;
		10'd841: data = 2'd1;
		10'd842: data = 2'd1;
		10'd843: data = 2'd2;
		10'd844: data = 2'd0;
		10'd845: data = 2'd1;
		10'd846: data = 2'd1;
		10'd847: data = 2'd3;
		10'd848: data = 2'd0;
		10'd849: data = 2'd1;
		10'd850: data = 2'd1;
		10'd851: data = 2'd3;
		10'd852: data = 2'd0;
		10'd853: data = 2'd0;
		10'd854: data = 2'd1;
		10'd855: data = 2'd3;
		10'd856: data = 2'd0;
		10'd857: data = 2'd0;
		10'd858: data = 2'd2;
		10'd859: data = 2'd3;
		10'd860: data = 2'd0;
		10'd861: data = 2'd0;
		10'd862: data = 2'd2;
		10'd863: data = 2'd3;
		10'd864: data = 2'd0;
		10'd865: data = 2'd0;
		10'd866: data = 2'd2;
		10'd867: data = 2'd3;
		10'd868: data = 2'd0;
		10'd869: data = 2'd0;
		10'd870: data = 2'd0;
		10'd871: data = 2'd3;
		10'd872: data = 2'd0;
		10'd873: data = 2'd0;
		10'd874: data = 2'd1;
		10'd875: data = 2'd3;
		10'd876: data = 2'd0;
		10'd877: data = 2'd0;
		10'd878: data = 2'd1;
		10'd879: data = 2'd3;
		10'd880: data = 2'd0;
		10'd881: data = 2'd0;
		10'd882: data = 2'd0;
		10'd883: data = 2'd3;
		10'd884: data = 2'd0;
		10'd885: data = 2'd1;
		10'd886: data = 2'd0;
		10'd887: data = 2'd3;
		10'd888: data = 2'd0;
		10'd889: data = 2'd1;
		10'd890: data = 2'd0;
		10'd891: data = 2'd2;
		10'd892: data = 2'd0;
		10'd893: data = 2'd1;
		10'd894: data = 2'd1;
		10'd895: data = 2'd1;
		10'd896: data = 2'd0;
		10'd897: data = 2'd1;
		10'd898: data = 2'd1;
		10'd899: data = 2'd1;
		10'd900: data = 2'd0;
		10'd901: data = 2'd1;
		10'd902: data = 2'd2;
		10'd903: data = 2'd2;
		10'd904: data = 2'd0;
		10'd905: data = 2'd1;
		10'd906: data = 2'd1;
		10'd907: data = 2'd3;
		10'd908: data = 2'd0;
		10'd909: data = 2'd1;
		10'd910: data = 2'd1;
		10'd911: data = 2'd3;
		10'd912: data = 2'd0;
		10'd913: data = 2'd1;
		10'd914: data = 2'd1;
		10'd915: data = 2'd3;
		10'd916: data = 2'd0;
		10'd917: data = 2'd0;
		10'd918: data = 2'd2;
		10'd919: data = 2'd3;
		10'd920: data = 2'd0;
		10'd921: data = 2'd0;
		10'd922: data = 2'd3;
		10'd923: data = 2'd3;
		10'd924: data = 2'd0;
		10'd925: data = 2'd0;
		10'd926: data = 2'd3;
		10'd927: data = 2'd3;
		10'd928: data = 2'd0;
		10'd929: data = 2'd0;
		10'd930: data = 2'd3;
		10'd931: data = 2'd3;
		10'd932: data = 2'd0;
		10'd933: data = 2'd0;
		10'd934: data = 2'd2;
		10'd935: data = 2'd3;
		10'd936: data = 2'd0;
		10'd937: data = 2'd0;
		10'd938: data = 2'd0;
		10'd939: data = 2'd3;
		10'd940: data = 2'd0;
		10'd941: data = 2'd0;
		10'd942: data = 2'd1;
		10'd943: data = 2'd3;
		10'd944: data = 2'd0;
		10'd945: data = 2'd0;
		10'd946: data = 2'd1;
		10'd947: data = 2'd3;
		10'd948: data = 2'd0;
		10'd949: data = 2'd0;
		10'd950: data = 2'd0;
		10'd951: data = 2'd3;
		10'd952: data = 2'd0;
		10'd953: data = 2'd1;
		10'd954: data = 2'd0;
		10'd955: data = 2'd3;
		10'd956: data = 2'd0;
		10'd957: data = 2'd1;
		10'd958: data = 2'd0;
		10'd959: data = 2'd2;
		10'd960: data = 2'd0;
		10'd961: data = 2'd1;
		10'd962: data = 2'd0;
		10'd963: data = 2'd2;
		10'd964: data = 2'd0;
		10'd965: data = 2'd1;
		10'd966: data = 2'd2;
		10'd967: data = 2'd2;
		10'd968: data = 2'd0;
		10'd969: data = 2'd1;
		10'd970: data = 2'd1;
		10'd971: data = 2'd2;
		10'd972: data = 2'd0;
		10'd973: data = 2'd1;
		10'd974: data = 2'd0;
		10'd975: data = 2'd3;
		10'd976: data = 2'd0;
		10'd977: data = 2'd0;
		10'd978: data = 2'd2;
		10'd979: data = 2'd3;
		10'd980: data = 2'd0;
		10'd981: data = 2'd0;
		10'd982: data = 2'd2;
		10'd983: data = 2'd3;
		10'd984: data = 2'd0;
		10'd985: data = 2'd0;
		10'd986: data = 2'd3;
		10'd987: data = 2'd3;
		10'd988: data = 2'd0;
		10'd989: data = 2'd0;
		10'd990: data = 2'd3;
		10'd991: data = 2'd3;
		10'd992: data = 2'd0;
		10'd993: data = 2'd0;
		10'd994: data = 2'd3;
		10'd995: data = 2'd3;
		10'd996: data = 2'd0;
		10'd997: data = 2'd0;
		10'd998: data = 2'd3;
		10'd999: data = 2'd3;
		10'd1000: data = 2'd0;
		10'd1001: data = 2'd0;
		10'd1002: data = 2'd2;
		10'd1003: data = 2'd3;
		10'd1004: data = 2'd0;
		10'd1005: data = 2'd0;
		10'd1006: data = 2'd2;
		10'd1007: data = 2'd3;
		10'd1008: data = 2'd0;
		10'd1009: data = 2'd0;
		10'd1010: data = 2'd1;
		10'd1011: data = 2'd3;
		10'd1012: data = 2'd0;
		10'd1013: data = 2'd0;
		10'd1014: data = 2'd1;
		10'd1015: data = 2'd3;
		10'd1016: data = 2'd0;
		10'd1017: data = 2'd0;
		10'd1018: data = 2'd0;
		10'd1019: data = 2'd3;
		10'd1020: data = 2'd0;
		10'd1021: data = 2'd1;
		10'd1022: data = 2'd0;
		10'd1023: data = 2'd3;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N0(address, data);
input wire [11:0] address;
output reg [3:0] data;

wire [4:0] i; layer1_N0_idx_1 idx_1_inst(address[11:2], i);
wire [1:0] t; layer1_N0_rsh_1 rsh_1_inst(address[11:2], t);
wire [3:0] b; layer1_N0_2 layer1_N0_2_inst(address[11:2], b);
wire [2:0] u; layer1_N0_ust_1 ust_1_inst({i, address[1:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule
