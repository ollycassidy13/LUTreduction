
module layer0_N23_ust_3(address, data);
input wire [5:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		6'd0: data = 2'd0;
		6'd1: data = 2'd0;
		6'd2: data = 2'd0;
		6'd3: data = 2'd1;
		6'd4: data = 2'd1;
		6'd5: data = 2'd2;
		6'd6: data = 2'd2;
		6'd7: data = 2'd3;
		6'd8: data = 2'd0;
		6'd9: data = 2'd0;
		6'd10: data = 2'd0;
		6'd11: data = 2'd0;
		6'd12: data = 2'd1;
		6'd13: data = 2'd1;
		6'd14: data = 2'd2;
		6'd15: data = 2'd3;
		6'd16: data = 2'd0;
		6'd17: data = 2'd0;
		6'd18: data = 2'd1;
		6'd19: data = 2'd1;
		6'd20: data = 2'd1;
		6'd21: data = 2'd2;
		6'd22: data = 2'd3;
		6'd23: data = 2'd3;
		6'd24: data = 2'd0;
		6'd25: data = 2'd0;
		6'd26: data = 2'd1;
		6'd27: data = 2'd1;
		6'd28: data = 2'd2;
		6'd29: data = 2'd2;
		6'd30: data = 2'd3;
		6'd31: data = 2'd3;
		6'd32: data = 2'd0;
		6'd33: data = 2'd0;
		6'd34: data = 2'd1;
		6'd35: data = 2'd1;
		6'd36: data = 2'd1;
		6'd37: data = 2'd2;
		6'd38: data = 2'd2;
		6'd39: data = 2'd3;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N23_idx_3(address, data);
input wire [3:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		4'd0: data = 3'd1;
		4'd1: data = 3'd1;
		4'd2: data = 3'd1;
		4'd3: data = 3'd0;
		4'd4: data = 3'd0;
		4'd5: data = 3'd0;
		4'd6: data = 3'd0;
		4'd7: data = 3'd0;
		4'd8: data = 3'd0;
		4'd9: data = 3'd4;
		4'd10: data = 3'd2;
		4'd11: data = 3'd2;
		4'd12: data = 3'd2;
		4'd13: data = 3'd3;
		4'd14: data = 3'd3;
		4'd15: data = 3'd3;
		default: data = 3'd0;
	endcase
end
endmodule

module layer0_N23_lb_3(address, data);
input wire [6:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		7'd0: data = 2'd2;
		7'd1: data = 2'd2;
		7'd2: data = 2'd2;
		7'd3: data = 2'd2;
		7'd4: data = 2'd0;
		7'd5: data = 2'd2;
		7'd6: data = 2'd1;
		7'd7: data = 2'd0;
		7'd8: data = 2'd2;
		7'd9: data = 2'd3;
		7'd10: data = 2'd3;
		7'd11: data = 2'd3;
		7'd12: data = 2'd0;
		7'd13: data = 2'd3;
		7'd14: data = 2'd1;
		7'd15: data = 2'd0;
		7'd16: data = 2'd3;
		7'd17: data = 2'd3;
		7'd18: data = 2'd3;
		7'd19: data = 2'd3;
		7'd20: data = 2'd1;
		7'd21: data = 2'd3;
		7'd22: data = 2'd2;
		7'd23: data = 2'd1;
		7'd24: data = 2'd3;
		7'd25: data = 2'd3;
		7'd26: data = 2'd3;
		7'd27: data = 2'd0;
		7'd28: data = 2'd2;
		7'd29: data = 2'd0;
		7'd30: data = 2'd2;
		7'd31: data = 2'd1;
		7'd32: data = 2'd3;
		7'd33: data = 2'd3;
		7'd34: data = 2'd3;
		7'd35: data = 2'd0;
		7'd36: data = 2'd2;
		7'd37: data = 2'd0;
		7'd38: data = 2'd2;
		7'd39: data = 2'd1;
		7'd40: data = 2'd3;
		7'd41: data = 2'd3;
		7'd42: data = 2'd3;
		7'd43: data = 2'd1;
		7'd44: data = 2'd2;
		7'd45: data = 2'd0;
		7'd46: data = 2'd3;
		7'd47: data = 2'd2;
		7'd48: data = 2'd3;
		7'd49: data = 2'd3;
		7'd50: data = 2'd3;
		7'd51: data = 2'd1;
		7'd52: data = 2'd2;
		7'd53: data = 2'd1;
		7'd54: data = 2'd3;
		7'd55: data = 2'd2;
		7'd56: data = 2'd2;
		7'd57: data = 2'd3;
		7'd58: data = 2'd3;
		7'd59: data = 2'd1;
		7'd60: data = 2'd3;
		7'd61: data = 2'd1;
		7'd62: data = 2'd3;
		7'd63: data = 2'd2;
		7'd64: data = 2'd2;
		7'd65: data = 2'd3;
		7'd66: data = 2'd3;
		7'd67: data = 2'd1;
		7'd68: data = 2'd3;
		7'd69: data = 2'd1;
		7'd70: data = 2'd3;
		7'd71: data = 2'd2;
		7'd72: data = 2'd2;
		7'd73: data = 2'd3;
		7'd74: data = 2'd0;
		7'd75: data = 2'd1;
		7'd76: data = 2'd3;
		7'd77: data = 2'd1;
		7'd78: data = 2'd3;
		7'd79: data = 2'd3;
		7'd80: data = 2'd1;
		7'd81: data = 2'd3;
		7'd82: data = 2'd0;
		7'd83: data = 2'd1;
		7'd84: data = 2'd3;
		7'd85: data = 2'd1;
		7'd86: data = 2'd0;
		7'd87: data = 2'd3;
		7'd88: data = 2'd1;
		7'd89: data = 2'd2;
		7'd90: data = 2'd0;
		7'd91: data = 2'd2;
		7'd92: data = 2'd3;
		7'd93: data = 2'd1;
		7'd94: data = 2'd0;
		7'd95: data = 2'd3;
		7'd96: data = 2'd0;
		7'd97: data = 2'd2;
		7'd98: data = 2'd0;
		7'd99: data = 2'd2;
		7'd100: data = 2'd3;
		7'd101: data = 2'd2;
		7'd102: data = 2'd0;
		7'd103: data = 2'd3;
		7'd104: data = 2'd0;
		7'd105: data = 2'd2;
		7'd106: data = 2'd0;
		7'd107: data = 2'd2;
		7'd108: data = 2'd0;
		7'd109: data = 2'd2;
		7'd110: data = 2'd0;
		7'd111: data = 2'd3;
		7'd112: data = 2'd0;
		7'd113: data = 2'd2;
		7'd114: data = 2'd0;
		7'd115: data = 2'd2;
		7'd116: data = 2'd0;
		7'd117: data = 2'd2;
		7'd118: data = 2'd1;
		7'd119: data = 2'd3;
		7'd120: data = 2'd0;
		7'd121: data = 2'd2;
		7'd122: data = 2'd0;
		7'd123: data = 2'd2;
		7'd124: data = 2'd0;
		7'd125: data = 2'd2;
		7'd126: data = 2'd1;
		7'd127: data = 2'd3;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N23_3(address, data);
input wire [6:0] address;
output reg [3:0] data;

wire [2:0] i; layer0_N23_idx_3 idx_3_inst(address[6:3], i);
wire [1:0] lb; layer0_N23_lb_3 lb_3_inst(address, lb);
wire [1:0] u; layer0_N23_ust_3 ust_3_inst({i, address[2:0]}, u);

always @(*) begin
	data = {u, lb};
end
endmodule

module layer0_N23_ust_2(address, data);
input wire [5:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		6'd0: data = 2'd1;
		6'd1: data = 2'd0;
		6'd2: data = 2'd2;
		6'd3: data = 2'd1;
		6'd4: data = 2'd1;
		6'd5: data = 2'd0;
		6'd6: data = 2'd2;
		6'd7: data = 2'd2;
		6'd8: data = 2'd2;
		6'd9: data = 2'd0;
		6'd10: data = 2'd3;
		6'd11: data = 2'd1;
		6'd12: data = 2'd0;
		6'd13: data = 2'd0;
		6'd14: data = 2'd2;
		6'd15: data = 2'd1;
		6'd16: data = 2'd2;
		6'd17: data = 2'd0;
		6'd18: data = 2'd3;
		6'd19: data = 2'd2;
		6'd20: data = 2'd1;
		6'd21: data = 2'd0;
		6'd22: data = 2'd3;
		6'd23: data = 2'd2;
		6'd24: data = 2'd0;
		6'd25: data = 2'd0;
		6'd26: data = 2'd2;
		6'd27: data = 2'd2;
		6'd28: data = 2'd2;
		6'd29: data = 2'd0;
		6'd30: data = 2'd2;
		6'd31: data = 2'd0;
		6'd32: data = 2'd1;
		6'd33: data = 2'd0;
		6'd34: data = 2'd2;
		6'd35: data = 2'd0;
		6'd36: data = 2'd2;
		6'd37: data = 2'd0;
		6'd38: data = 2'd2;
		6'd39: data = 2'd1;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N23_idx_2(address, data);
input wire [6:0] address;
output reg [3:0] data;

always @(*) begin
	case(address)
		7'd0: data = 4'd2;
		7'd1: data = 4'd8;
		7'd2: data = 4'd7;
		7'd3: data = 4'd2;
		7'd4: data = 4'd2;
		7'd5: data = 4'd4;
		7'd6: data = 4'd0;
		7'd7: data = 4'd5;
		7'd8: data = 4'd2;
		7'd9: data = 4'd0;
		7'd10: data = 4'd2;
		7'd11: data = 4'd7;
		7'd12: data = 4'd4;
		7'd13: data = 4'd0;
		7'd14: data = 4'd1;
		7'd15: data = 4'd5;
		7'd16: data = 4'd0;
		7'd17: data = 4'd0;
		7'd18: data = 4'd2;
		7'd19: data = 4'd2;
		7'd20: data = 4'd9;
		7'd21: data = 4'd0;
		7'd22: data = 4'd3;
		7'd23: data = 4'd6;
		7'd24: data = 4'd0;
		7'd25: data = 4'd0;
		7'd26: data = 4'd2;
		7'd27: data = 4'd0;
		7'd28: data = 4'd0;
		7'd29: data = 4'd0;
		7'd30: data = 4'd3;
		7'd31: data = 4'd1;
		7'd32: data = 4'd0;
		7'd33: data = 4'd0;
		7'd34: data = 4'd2;
		7'd35: data = 4'd0;
		7'd36: data = 4'd0;
		7'd37: data = 4'd0;
		7'd38: data = 4'd1;
		7'd39: data = 4'd1;
		7'd40: data = 4'd0;
		7'd41: data = 4'd0;
		7'd42: data = 4'd0;
		7'd43: data = 4'd0;
		7'd44: data = 4'd0;
		7'd45: data = 4'd0;
		7'd46: data = 4'd1;
		7'd47: data = 4'd1;
		7'd48: data = 4'd0;
		7'd49: data = 4'd0;
		7'd50: data = 4'd0;
		7'd51: data = 4'd1;
		7'd52: data = 4'd0;
		7'd53: data = 4'd1;
		7'd54: data = 4'd3;
		7'd55: data = 4'd4;
		7'd56: data = 4'd1;
		7'd57: data = 4'd0;
		7'd58: data = 4'd0;
		7'd59: data = 4'd0;
		7'd60: data = 4'd1;
		7'd61: data = 4'd1;
		7'd62: data = 4'd3;
		7'd63: data = 4'd4;
		7'd64: data = 4'd0;
		7'd65: data = 4'd0;
		7'd66: data = 4'd0;
		7'd67: data = 4'd0;
		7'd68: data = 4'd0;
		7'd69: data = 4'd1;
		7'd70: data = 4'd6;
		7'd71: data = 4'd4;
		7'd72: data = 4'd0;
		7'd73: data = 4'd0;
		7'd74: data = 4'd0;
		7'd75: data = 4'd0;
		7'd76: data = 4'd0;
		7'd77: data = 4'd0;
		7'd78: data = 4'd1;
		7'd79: data = 4'd0;
		7'd80: data = 4'd1;
		7'd81: data = 4'd0;
		7'd82: data = 4'd1;
		7'd83: data = 4'd0;
		7'd84: data = 4'd0;
		7'd85: data = 4'd0;
		7'd86: data = 4'd3;
		7'd87: data = 4'd0;
		7'd88: data = 4'd1;
		7'd89: data = 4'd0;
		7'd90: data = 4'd1;
		7'd91: data = 4'd0;
		7'd92: data = 4'd0;
		7'd93: data = 4'd1;
		7'd94: data = 4'd3;
		7'd95: data = 4'd0;
		7'd96: data = 4'd1;
		7'd97: data = 4'd0;
		7'd98: data = 4'd0;
		7'd99: data = 4'd1;
		7'd100: data = 4'd0;
		7'd101: data = 4'd1;
		7'd102: data = 4'd6;
		7'd103: data = 4'd0;
		7'd104: data = 4'd1;
		7'd105: data = 4'd0;
		7'd106: data = 4'd0;
		7'd107: data = 4'd0;
		7'd108: data = 4'd1;
		7'd109: data = 4'd1;
		7'd110: data = 4'd5;
		7'd111: data = 4'd0;
		7'd112: data = 4'd0;
		7'd113: data = 4'd0;
		7'd114: data = 4'd0;
		7'd115: data = 4'd0;
		7'd116: data = 4'd0;
		7'd117: data = 4'd1;
		7'd118: data = 4'd3;
		7'd119: data = 4'd0;
		7'd120: data = 4'd0;
		7'd121: data = 4'd0;
		7'd122: data = 4'd0;
		7'd123: data = 4'd0;
		7'd124: data = 4'd0;
		7'd125: data = 4'd1;
		7'd126: data = 4'd3;
		7'd127: data = 4'd0;
		default: data = 4'd0;
	endcase
end
endmodule

module layer0_N23_rsh_2(address, data);
input wire [6:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		7'd0: data = 2'd1;
		7'd1: data = 2'd0;
		7'd2: data = 2'd0;
		7'd3: data = 2'd0;
		7'd4: data = 2'd0;
		7'd5: data = 2'd0;
		7'd6: data = 2'd0;
		7'd7: data = 2'd0;
		7'd8: data = 2'd1;
		7'd9: data = 2'd1;
		7'd10: data = 2'd1;
		7'd11: data = 2'd0;
		7'd12: data = 2'd0;
		7'd13: data = 2'd0;
		7'd14: data = 2'd0;
		7'd15: data = 2'd0;
		7'd16: data = 2'd2;
		7'd17: data = 2'd2;
		7'd18: data = 2'd1;
		7'd19: data = 2'd0;
		7'd20: data = 2'd0;
		7'd21: data = 2'd0;
		7'd22: data = 2'd0;
		7'd23: data = 2'd0;
		7'd24: data = 2'd2;
		7'd25: data = 2'd2;
		7'd26: data = 2'd1;
		7'd27: data = 2'd0;
		7'd28: data = 2'd0;
		7'd29: data = 2'd0;
		7'd30: data = 2'd0;
		7'd31: data = 2'd0;
		7'd32: data = 2'd2;
		7'd33: data = 2'd2;
		7'd34: data = 2'd1;
		7'd35: data = 2'd0;
		7'd36: data = 2'd0;
		7'd37: data = 2'd0;
		7'd38: data = 2'd0;
		7'd39: data = 2'd0;
		7'd40: data = 2'd2;
		7'd41: data = 2'd2;
		7'd42: data = 2'd0;
		7'd43: data = 2'd1;
		7'd44: data = 2'd0;
		7'd45: data = 2'd0;
		7'd46: data = 2'd1;
		7'd47: data = 2'd1;
		7'd48: data = 2'd2;
		7'd49: data = 2'd2;
		7'd50: data = 2'd0;
		7'd51: data = 2'd1;
		7'd52: data = 2'd0;
		7'd53: data = 2'd1;
		7'd54: data = 2'd0;
		7'd55: data = 2'd1;
		7'd56: data = 2'd1;
		7'd57: data = 2'd2;
		7'd58: data = 2'd0;
		7'd59: data = 2'd0;
		7'd60: data = 2'd1;
		7'd61: data = 2'd1;
		7'd62: data = 2'd0;
		7'd63: data = 2'd1;
		7'd64: data = 2'd1;
		7'd65: data = 2'd2;
		7'd66: data = 2'd0;
		7'd67: data = 2'd0;
		7'd68: data = 2'd0;
		7'd69: data = 2'd1;
		7'd70: data = 2'd0;
		7'd71: data = 2'd1;
		7'd72: data = 2'd2;
		7'd73: data = 2'd2;
		7'd74: data = 2'd1;
		7'd75: data = 2'd0;
		7'd76: data = 2'd0;
		7'd77: data = 2'd0;
		7'd78: data = 2'd0;
		7'd79: data = 2'd2;
		7'd80: data = 2'd1;
		7'd81: data = 2'd2;
		7'd82: data = 2'd1;
		7'd83: data = 2'd0;
		7'd84: data = 2'd0;
		7'd85: data = 2'd0;
		7'd86: data = 2'd0;
		7'd87: data = 2'd2;
		7'd88: data = 2'd1;
		7'd89: data = 2'd0;
		7'd90: data = 2'd1;
		7'd91: data = 2'd1;
		7'd92: data = 2'd0;
		7'd93: data = 2'd0;
		7'd94: data = 2'd0;
		7'd95: data = 2'd2;
		7'd96: data = 2'd1;
		7'd97: data = 2'd0;
		7'd98: data = 2'd0;
		7'd99: data = 2'd1;
		7'd100: data = 2'd0;
		7'd101: data = 2'd1;
		7'd102: data = 2'd0;
		7'd103: data = 2'd2;
		7'd104: data = 2'd1;
		7'd105: data = 2'd0;
		7'd106: data = 2'd0;
		7'd107: data = 2'd0;
		7'd108: data = 2'd1;
		7'd109: data = 2'd1;
		7'd110: data = 2'd0;
		7'd111: data = 2'd2;
		7'd112: data = 2'd1;
		7'd113: data = 2'd0;
		7'd114: data = 2'd0;
		7'd115: data = 2'd0;
		7'd116: data = 2'd0;
		7'd117: data = 2'd1;
		7'd118: data = 2'd0;
		7'd119: data = 2'd2;
		7'd120: data = 2'd1;
		7'd121: data = 2'd0;
		7'd122: data = 2'd0;
		7'd123: data = 2'd0;
		7'd124: data = 2'd0;
		7'd125: data = 2'd0;
		7'd126: data = 2'd0;
		7'd127: data = 2'd2;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N23_2(address, data);
input wire [8:0] address;
output reg [3:0] data;

wire [3:0] i; layer0_N23_idx_2 idx_2_inst(address[8:2], i);
wire [1:0] t; layer0_N23_rsh_2 rsh_2_inst(address[8:2], t);
wire [3:0] b; layer0_N23_3 layer0_N23_3_inst(address[8:2], b);
wire [1:0] u; layer0_N23_ust_2 ust_2_inst({i, address[1:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule

module layer0_N23_ust_1(address, data);
input wire [8:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		9'd0: data = 3'd4;
		9'd1: data = 3'd3;
		9'd2: data = 3'd3;
		9'd3: data = 3'd2;
		9'd4: data = 3'd1;
		9'd5: data = 3'd1;
		9'd6: data = 3'd1;
		9'd7: data = 3'd0;
		9'd8: data = 3'd2;
		9'd9: data = 3'd2;
		9'd10: data = 3'd1;
		9'd11: data = 3'd1;
		9'd12: data = 3'd1;
		9'd13: data = 3'd0;
		9'd14: data = 3'd0;
		9'd15: data = 3'd0;
		9'd16: data = 3'd2;
		9'd17: data = 3'd2;
		9'd18: data = 3'd2;
		9'd19: data = 3'd1;
		9'd20: data = 3'd1;
		9'd21: data = 3'd1;
		9'd22: data = 3'd0;
		9'd23: data = 3'd0;
		9'd24: data = 3'd2;
		9'd25: data = 3'd2;
		9'd26: data = 3'd2;
		9'd27: data = 3'd2;
		9'd28: data = 3'd1;
		9'd29: data = 3'd1;
		9'd30: data = 3'd1;
		9'd31: data = 3'd0;
		9'd32: data = 3'd2;
		9'd33: data = 3'd2;
		9'd34: data = 3'd2;
		9'd35: data = 3'd2;
		9'd36: data = 3'd2;
		9'd37: data = 3'd1;
		9'd38: data = 3'd1;
		9'd39: data = 3'd0;
		9'd40: data = 3'd1;
		9'd41: data = 3'd1;
		9'd42: data = 3'd1;
		9'd43: data = 3'd1;
		9'd44: data = 3'd1;
		9'd45: data = 3'd1;
		9'd46: data = 3'd1;
		9'd47: data = 3'd0;
		9'd48: data = 3'd1;
		9'd49: data = 3'd1;
		9'd50: data = 3'd1;
		9'd51: data = 3'd1;
		9'd52: data = 3'd1;
		9'd53: data = 3'd1;
		9'd54: data = 3'd0;
		9'd55: data = 3'd0;
		9'd56: data = 3'd2;
		9'd57: data = 3'd1;
		9'd58: data = 3'd1;
		9'd59: data = 3'd0;
		9'd60: data = 3'd0;
		9'd61: data = 3'd0;
		9'd62: data = 3'd0;
		9'd63: data = 3'd0;
		9'd64: data = 3'd2;
		9'd65: data = 3'd2;
		9'd66: data = 3'd1;
		9'd67: data = 3'd1;
		9'd68: data = 3'd1;
		9'd69: data = 3'd1;
		9'd70: data = 3'd1;
		9'd71: data = 3'd0;
		9'd72: data = 3'd2;
		9'd73: data = 3'd2;
		9'd74: data = 3'd1;
		9'd75: data = 3'd1;
		9'd76: data = 3'd1;
		9'd77: data = 3'd1;
		9'd78: data = 3'd0;
		9'd79: data = 3'd0;
		9'd80: data = 3'd2;
		9'd81: data = 3'd1;
		9'd82: data = 3'd1;
		9'd83: data = 3'd1;
		9'd84: data = 3'd1;
		9'd85: data = 3'd1;
		9'd86: data = 3'd1;
		9'd87: data = 3'd0;
		9'd88: data = 3'd2;
		9'd89: data = 3'd2;
		9'd90: data = 3'd1;
		9'd91: data = 3'd1;
		9'd92: data = 3'd0;
		9'd93: data = 3'd0;
		9'd94: data = 3'd0;
		9'd95: data = 3'd0;
		9'd96: data = 3'd2;
		9'd97: data = 3'd2;
		9'd98: data = 3'd2;
		9'd99: data = 3'd1;
		9'd100: data = 3'd1;
		9'd101: data = 3'd0;
		9'd102: data = 3'd0;
		9'd103: data = 3'd0;
		9'd104: data = 3'd2;
		9'd105: data = 3'd1;
		9'd106: data = 3'd1;
		9'd107: data = 3'd1;
		9'd108: data = 3'd1;
		9'd109: data = 3'd0;
		9'd110: data = 3'd0;
		9'd111: data = 3'd0;
		9'd112: data = 3'd2;
		9'd113: data = 3'd2;
		9'd114: data = 3'd2;
		9'd115: data = 3'd1;
		9'd116: data = 3'd1;
		9'd117: data = 3'd1;
		9'd118: data = 3'd1;
		9'd119: data = 3'd0;
		9'd120: data = 3'd3;
		9'd121: data = 3'd2;
		9'd122: data = 3'd2;
		9'd123: data = 3'd1;
		9'd124: data = 3'd1;
		9'd125: data = 3'd1;
		9'd126: data = 3'd0;
		9'd127: data = 3'd0;
		9'd128: data = 3'd2;
		9'd129: data = 3'd1;
		9'd130: data = 3'd1;
		9'd131: data = 3'd1;
		9'd132: data = 3'd1;
		9'd133: data = 3'd1;
		9'd134: data = 3'd0;
		9'd135: data = 3'd0;
		9'd136: data = 3'd0;
		9'd137: data = 3'd0;
		9'd138: data = 3'd0;
		9'd139: data = 3'd0;
		9'd140: data = 3'd0;
		9'd141: data = 3'd0;
		9'd142: data = 3'd0;
		9'd143: data = 3'd1;
		9'd144: data = 3'd3;
		9'd145: data = 3'd2;
		9'd146: data = 3'd2;
		9'd147: data = 3'd1;
		9'd148: data = 3'd1;
		9'd149: data = 3'd1;
		9'd150: data = 3'd1;
		9'd151: data = 3'd0;
		9'd152: data = 3'd3;
		9'd153: data = 3'd2;
		9'd154: data = 3'd2;
		9'd155: data = 3'd2;
		9'd156: data = 3'd1;
		9'd157: data = 3'd1;
		9'd158: data = 3'd1;
		9'd159: data = 3'd0;
		9'd160: data = 3'd2;
		9'd161: data = 3'd2;
		9'd162: data = 3'd2;
		9'd163: data = 3'd2;
		9'd164: data = 3'd1;
		9'd165: data = 3'd1;
		9'd166: data = 3'd0;
		9'd167: data = 3'd0;
		9'd168: data = 3'd3;
		9'd169: data = 3'd3;
		9'd170: data = 3'd2;
		9'd171: data = 3'd1;
		9'd172: data = 3'd1;
		9'd173: data = 3'd1;
		9'd174: data = 3'd0;
		9'd175: data = 3'd0;
		9'd176: data = 3'd3;
		9'd177: data = 3'd3;
		9'd178: data = 3'd2;
		9'd179: data = 3'd1;
		9'd180: data = 3'd1;
		9'd181: data = 3'd0;
		9'd182: data = 3'd0;
		9'd183: data = 3'd0;
		9'd184: data = 3'd1;
		9'd185: data = 3'd1;
		9'd186: data = 3'd1;
		9'd187: data = 3'd0;
		9'd188: data = 3'd0;
		9'd189: data = 3'd0;
		9'd190: data = 3'd0;
		9'd191: data = 3'd1;
		9'd192: data = 3'd3;
		9'd193: data = 3'd2;
		9'd194: data = 3'd1;
		9'd195: data = 3'd1;
		9'd196: data = 3'd1;
		9'd197: data = 3'd1;
		9'd198: data = 3'd0;
		9'd199: data = 3'd0;
		9'd200: data = 3'd0;
		9'd201: data = 3'd0;
		9'd202: data = 3'd0;
		9'd203: data = 3'd0;
		9'd204: data = 3'd0;
		9'd205: data = 3'd0;
		9'd206: data = 3'd1;
		9'd207: data = 3'd1;
		9'd208: data = 3'd0;
		9'd209: data = 3'd0;
		9'd210: data = 3'd1;
		9'd211: data = 3'd1;
		9'd212: data = 3'd1;
		9'd213: data = 3'd1;
		9'd214: data = 3'd1;
		9'd215: data = 3'd1;
		9'd216: data = 3'd0;
		9'd217: data = 3'd0;
		9'd218: data = 3'd0;
		9'd219: data = 3'd0;
		9'd220: data = 3'd0;
		9'd221: data = 3'd1;
		9'd222: data = 3'd1;
		9'd223: data = 3'd1;
		9'd224: data = 3'd3;
		9'd225: data = 3'd2;
		9'd226: data = 3'd2;
		9'd227: data = 3'd1;
		9'd228: data = 3'd1;
		9'd229: data = 3'd0;
		9'd230: data = 3'd0;
		9'd231: data = 3'd0;
		9'd232: data = 3'd2;
		9'd233: data = 3'd2;
		9'd234: data = 3'd2;
		9'd235: data = 3'd2;
		9'd236: data = 3'd1;
		9'd237: data = 3'd0;
		9'd238: data = 3'd0;
		9'd239: data = 3'd0;
		9'd240: data = 3'd2;
		9'd241: data = 3'd2;
		9'd242: data = 3'd2;
		9'd243: data = 3'd2;
		9'd244: data = 3'd2;
		9'd245: data = 3'd1;
		9'd246: data = 3'd0;
		9'd247: data = 3'd0;
		9'd248: data = 3'd3;
		9'd249: data = 3'd3;
		9'd250: data = 3'd2;
		9'd251: data = 3'd1;
		9'd252: data = 3'd1;
		9'd253: data = 3'd1;
		9'd254: data = 3'd1;
		9'd255: data = 3'd0;
		9'd256: data = 3'd1;
		9'd257: data = 3'd1;
		9'd258: data = 3'd0;
		9'd259: data = 3'd0;
		9'd260: data = 3'd0;
		9'd261: data = 3'd0;
		9'd262: data = 3'd0;
		9'd263: data = 3'd1;
		9'd264: data = 3'd1;
		9'd265: data = 3'd0;
		9'd266: data = 3'd0;
		9'd267: data = 3'd0;
		9'd268: data = 3'd0;
		9'd269: data = 3'd0;
		9'd270: data = 3'd0;
		9'd271: data = 3'd1;
		9'd272: data = 3'd3;
		9'd273: data = 3'd2;
		9'd274: data = 3'd1;
		9'd275: data = 3'd1;
		9'd276: data = 3'd1;
		9'd277: data = 3'd0;
		9'd278: data = 3'd0;
		9'd279: data = 3'd0;
		9'd280: data = 3'd3;
		9'd281: data = 3'd3;
		9'd282: data = 3'd2;
		9'd283: data = 3'd2;
		9'd284: data = 3'd1;
		9'd285: data = 3'd1;
		9'd286: data = 3'd1;
		9'd287: data = 3'd0;
		9'd288: data = 3'd2;
		9'd289: data = 3'd2;
		9'd290: data = 3'd2;
		9'd291: data = 3'd1;
		9'd292: data = 3'd0;
		9'd293: data = 3'd0;
		9'd294: data = 3'd0;
		9'd295: data = 3'd0;
		9'd296: data = 3'd1;
		9'd297: data = 3'd1;
		9'd298: data = 3'd1;
		9'd299: data = 3'd0;
		9'd300: data = 3'd0;
		9'd301: data = 3'd1;
		9'd302: data = 3'd1;
		9'd303: data = 3'd1;
		9'd304: data = 3'd0;
		9'd305: data = 3'd0;
		9'd306: data = 3'd0;
		9'd307: data = 3'd1;
		9'd308: data = 3'd1;
		9'd309: data = 3'd1;
		9'd310: data = 3'd1;
		9'd311: data = 3'd1;
		9'd312: data = 3'd1;
		9'd313: data = 3'd1;
		9'd314: data = 3'd0;
		9'd315: data = 3'd0;
		9'd316: data = 3'd0;
		9'd317: data = 3'd0;
		9'd318: data = 3'd1;
		9'd319: data = 3'd1;
		9'd320: data = 3'd1;
		9'd321: data = 3'd1;
		9'd322: data = 3'd1;
		9'd323: data = 3'd1;
		9'd324: data = 3'd0;
		9'd325: data = 3'd0;
		9'd326: data = 3'd0;
		9'd327: data = 3'd1;
		9'd328: data = 3'd0;
		9'd329: data = 3'd1;
		9'd330: data = 3'd1;
		9'd331: data = 3'd1;
		9'd332: data = 3'd1;
		9'd333: data = 3'd1;
		9'd334: data = 3'd1;
		9'd335: data = 3'd1;
		9'd336: data = 3'd1;
		9'd337: data = 3'd1;
		9'd338: data = 3'd1;
		9'd339: data = 3'd1;
		9'd340: data = 3'd0;
		9'd341: data = 3'd1;
		9'd342: data = 3'd0;
		9'd343: data = 3'd0;
		9'd344: data = 3'd2;
		9'd345: data = 3'd1;
		9'd346: data = 3'd0;
		9'd347: data = 3'd0;
		9'd348: data = 3'd0;
		9'd349: data = 3'd0;
		9'd350: data = 3'd0;
		9'd351: data = 3'd0;
		default: data = 3'd0;
	endcase
end
endmodule

module layer0_N23_idx_1(address, data);
input wire [8:0] address;
output reg [5:0] data;

always @(*) begin
	case(address)
		9'd0: data = 6'd12;
		9'd1: data = 6'd6;
		9'd2: data = 6'd2;
		9'd3: data = 6'd5;
		9'd4: data = 6'd19;
		9'd5: data = 6'd5;
		9'd6: data = 6'd0;
		9'd7: data = 6'd5;
		9'd8: data = 6'd1;
		9'd9: data = 6'd8;
		9'd10: data = 6'd12;
		9'd11: data = 6'd14;
		9'd12: data = 6'd15;
		9'd13: data = 6'd3;
		9'd14: data = 6'd12;
		9'd15: data = 6'd2;
		9'd16: data = 6'd1;
		9'd17: data = 6'd20;
		9'd18: data = 6'd0;
		9'd19: data = 6'd3;
		9'd20: data = 6'd7;
		9'd21: data = 6'd14;
		9'd22: data = 6'd7;
		9'd23: data = 6'd1;
		9'd24: data = 6'd28;
		9'd25: data = 6'd1;
		9'd26: data = 6'd0;
		9'd27: data = 6'd2;
		9'd28: data = 6'd29;
		9'd29: data = 6'd1;
		9'd30: data = 6'd0;
		9'd31: data = 6'd2;
		9'd32: data = 6'd1;
		9'd33: data = 6'd5;
		9'd34: data = 6'd2;
		9'd35: data = 6'd5;
		9'd36: data = 6'd15;
		9'd37: data = 6'd0;
		9'd38: data = 6'd0;
		9'd39: data = 6'd0;
		9'd40: data = 6'd1;
		9'd41: data = 6'd1;
		9'd42: data = 6'd1;
		9'd43: data = 6'd2;
		9'd44: data = 6'd0;
		9'd45: data = 6'd3;
		9'd46: data = 6'd18;
		9'd47: data = 6'd3;
		9'd48: data = 6'd9;
		9'd49: data = 6'd4;
		9'd50: data = 6'd9;
		9'd51: data = 6'd6;
		9'd52: data = 6'd13;
		9'd53: data = 6'd4;
		9'd54: data = 6'd0;
		9'd55: data = 6'd3;
		9'd56: data = 6'd15;
		9'd57: data = 6'd3;
		9'd58: data = 6'd0;
		9'd59: data = 6'd0;
		9'd60: data = 6'd20;
		9'd61: data = 6'd6;
		9'd62: data = 6'd0;
		9'd63: data = 6'd5;
		9'd64: data = 6'd1;
		9'd65: data = 6'd0;
		9'd66: data = 6'd12;
		9'd67: data = 6'd0;
		9'd68: data = 6'd2;
		9'd69: data = 6'd0;
		9'd70: data = 6'd19;
		9'd71: data = 6'd0;
		9'd72: data = 6'd0;
		9'd73: data = 6'd2;
		9'd74: data = 6'd1;
		9'd75: data = 6'd3;
		9'd76: data = 6'd0;
		9'd77: data = 6'd13;
		9'd78: data = 6'd7;
		9'd79: data = 6'd16;
		9'd80: data = 6'd2;
		9'd81: data = 6'd6;
		9'd82: data = 6'd8;
		9'd83: data = 6'd5;
		9'd84: data = 6'd10;
		9'd85: data = 6'd5;
		9'd86: data = 6'd9;
		9'd87: data = 6'd6;
		9'd88: data = 6'd21;
		9'd89: data = 6'd0;
		9'd90: data = 6'd22;
		9'd91: data = 6'd0;
		9'd92: data = 6'd30;
		9'd93: data = 6'd0;
		9'd94: data = 6'd0;
		9'd95: data = 6'd0;
		9'd96: data = 6'd1;
		9'd97: data = 6'd0;
		9'd98: data = 6'd1;
		9'd99: data = 6'd0;
		9'd100: data = 6'd2;
		9'd101: data = 6'd0;
		9'd102: data = 6'd18;
		9'd103: data = 6'd0;
		9'd104: data = 6'd0;
		9'd105: data = 6'd1;
		9'd106: data = 6'd1;
		9'd107: data = 6'd3;
		9'd108: data = 6'd11;
		9'd109: data = 6'd2;
		9'd110: data = 6'd0;
		9'd111: data = 6'd1;
		9'd112: data = 6'd2;
		9'd113: data = 6'd1;
		9'd114: data = 6'd1;
		9'd115: data = 6'd0;
		9'd116: data = 6'd0;
		9'd117: data = 6'd0;
		9'd118: data = 6'd1;
		9'd119: data = 6'd0;
		9'd120: data = 6'd31;
		9'd121: data = 6'd0;
		9'd122: data = 6'd22;
		9'd123: data = 6'd32;
		9'd124: data = 6'd4;
		9'd125: data = 6'd2;
		9'd126: data = 6'd0;
		9'd127: data = 6'd0;
		9'd128: data = 6'd0;
		9'd129: data = 6'd0;
		9'd130: data = 6'd1;
		9'd131: data = 6'd0;
		9'd132: data = 6'd9;
		9'd133: data = 6'd0;
		9'd134: data = 6'd14;
		9'd135: data = 6'd0;
		9'd136: data = 6'd3;
		9'd137: data = 6'd1;
		9'd138: data = 6'd9;
		9'd139: data = 6'd3;
		9'd140: data = 6'd1;
		9'd141: data = 6'd4;
		9'd142: data = 6'd0;
		9'd143: data = 6'd3;
		9'd144: data = 6'd2;
		9'd145: data = 6'd2;
		9'd146: data = 6'd1;
		9'd147: data = 6'd2;
		9'd148: data = 6'd1;
		9'd149: data = 6'd1;
		9'd150: data = 6'd1;
		9'd151: data = 6'd0;
		9'd152: data = 6'd11;
		9'd153: data = 6'd33;
		9'd154: data = 6'd21;
		9'd155: data = 6'd0;
		9'd156: data = 6'd4;
		9'd157: data = 6'd5;
		9'd158: data = 6'd0;
		9'd159: data = 6'd0;
		9'd160: data = 6'd3;
		9'd161: data = 6'd0;
		9'd162: data = 6'd0;
		9'd163: data = 6'd0;
		9'd164: data = 6'd1;
		9'd165: data = 6'd0;
		9'd166: data = 6'd8;
		9'd167: data = 6'd0;
		9'd168: data = 6'd7;
		9'd169: data = 6'd1;
		9'd170: data = 6'd2;
		9'd171: data = 6'd0;
		9'd172: data = 6'd9;
		9'd173: data = 6'd0;
		9'd174: data = 6'd13;
		9'd175: data = 6'd6;
		9'd176: data = 6'd0;
		9'd177: data = 6'd4;
		9'd178: data = 6'd3;
		9'd179: data = 6'd4;
		9'd180: data = 6'd2;
		9'd181: data = 6'd3;
		9'd182: data = 6'd7;
		9'd183: data = 6'd23;
		9'd184: data = 6'd34;
		9'd185: data = 6'd0;
		9'd186: data = 6'd35;
		9'd187: data = 6'd0;
		9'd188: data = 6'd4;
		9'd189: data = 6'd0;
		9'd190: data = 6'd0;
		9'd191: data = 6'd0;
		9'd192: data = 6'd0;
		9'd193: data = 6'd0;
		9'd194: data = 6'd0;
		9'd195: data = 6'd0;
		9'd196: data = 6'd11;
		9'd197: data = 6'd0;
		9'd198: data = 6'd1;
		9'd199: data = 6'd0;
		9'd200: data = 6'd0;
		9'd201: data = 6'd0;
		9'd202: data = 6'd2;
		9'd203: data = 6'd0;
		9'd204: data = 6'd8;
		9'd205: data = 6'd0;
		9'd206: data = 6'd9;
		9'd207: data = 6'd0;
		9'd208: data = 6'd16;
		9'd209: data = 6'd5;
		9'd210: data = 6'd4;
		9'd211: data = 6'd5;
		9'd212: data = 6'd3;
		9'd213: data = 6'd0;
		9'd214: data = 6'd0;
		9'd215: data = 6'd0;
		9'd216: data = 6'd24;
		9'd217: data = 6'd0;
		9'd218: data = 6'd11;
		9'd219: data = 6'd25;
		9'd220: data = 6'd0;
		9'd221: data = 6'd0;
		9'd222: data = 6'd0;
		9'd223: data = 6'd0;
		9'd224: data = 6'd13;
		9'd225: data = 6'd26;
		9'd226: data = 6'd3;
		9'd227: data = 6'd0;
		9'd228: data = 6'd0;
		9'd229: data = 6'd0;
		9'd230: data = 6'd1;
		9'd231: data = 6'd0;
		9'd232: data = 6'd0;
		9'd233: data = 6'd1;
		9'd234: data = 6'd7;
		9'd235: data = 6'd0;
		9'd236: data = 6'd2;
		9'd237: data = 6'd0;
		9'd238: data = 6'd1;
		9'd239: data = 6'd0;
		9'd240: data = 6'd10;
		9'd241: data = 6'd0;
		9'd242: data = 6'd10;
		9'd243: data = 6'd0;
		9'd244: data = 6'd6;
		9'd245: data = 6'd0;
		9'd246: data = 6'd13;
		9'd247: data = 6'd0;
		9'd248: data = 6'd15;
		9'd249: data = 6'd17;
		9'd250: data = 6'd36;
		9'd251: data = 6'd37;
		9'd252: data = 6'd0;
		9'd253: data = 6'd3;
		9'd254: data = 6'd0;
		9'd255: data = 6'd0;
		9'd256: data = 6'd4;
		9'd257: data = 6'd25;
		9'd258: data = 6'd2;
		9'd259: data = 6'd38;
		9'd260: data = 6'd0;
		9'd261: data = 6'd0;
		9'd262: data = 6'd1;
		9'd263: data = 6'd0;
		9'd264: data = 6'd11;
		9'd265: data = 6'd23;
		9'd266: data = 6'd0;
		9'd267: data = 6'd2;
		9'd268: data = 6'd2;
		9'd269: data = 6'd1;
		9'd270: data = 6'd1;
		9'd271: data = 6'd0;
		9'd272: data = 6'd1;
		9'd273: data = 6'd0;
		9'd274: data = 6'd0;
		9'd275: data = 6'd0;
		9'd276: data = 6'd5;
		9'd277: data = 6'd0;
		9'd278: data = 6'd10;
		9'd279: data = 6'd0;
		9'd280: data = 6'd18;
		9'd281: data = 6'd17;
		9'd282: data = 6'd12;
		9'd283: data = 6'd0;
		9'd284: data = 6'd0;
		9'd285: data = 6'd5;
		9'd286: data = 6'd0;
		9'd287: data = 6'd0;
		9'd288: data = 6'd3;
		9'd289: data = 6'd0;
		9'd290: data = 6'd14;
		9'd291: data = 6'd0;
		9'd292: data = 6'd0;
		9'd293: data = 6'd0;
		9'd294: data = 6'd12;
		9'd295: data = 6'd0;
		9'd296: data = 6'd11;
		9'd297: data = 6'd0;
		9'd298: data = 6'd0;
		9'd299: data = 6'd3;
		9'd300: data = 6'd7;
		9'd301: data = 6'd2;
		9'd302: data = 6'd2;
		9'd303: data = 6'd2;
		9'd304: data = 6'd1;
		9'd305: data = 6'd1;
		9'd306: data = 6'd0;
		9'd307: data = 6'd0;
		9'd308: data = 6'd0;
		9'd309: data = 6'd0;
		9'd310: data = 6'd1;
		9'd311: data = 6'd0;
		9'd312: data = 6'd0;
		9'd313: data = 6'd27;
		9'd314: data = 6'd14;
		9'd315: data = 6'd0;
		9'd316: data = 6'd0;
		9'd317: data = 6'd0;
		9'd318: data = 6'd0;
		9'd319: data = 6'd0;
		9'd320: data = 6'd8;
		9'd321: data = 6'd26;
		9'd322: data = 6'd9;
		9'd323: data = 6'd0;
		9'd324: data = 6'd7;
		9'd325: data = 6'd0;
		9'd326: data = 6'd2;
		9'd327: data = 6'd0;
		9'd328: data = 6'd9;
		9'd329: data = 6'd0;
		9'd330: data = 6'd1;
		9'd331: data = 6'd0;
		9'd332: data = 6'd0;
		9'd333: data = 6'd4;
		9'd334: data = 6'd3;
		9'd335: data = 6'd3;
		9'd336: data = 6'd2;
		9'd337: data = 6'd3;
		9'd338: data = 6'd1;
		9'd339: data = 6'd2;
		9'd340: data = 6'd1;
		9'd341: data = 6'd1;
		9'd342: data = 6'd1;
		9'd343: data = 6'd39;
		9'd344: data = 6'd11;
		9'd345: data = 6'd0;
		9'd346: data = 6'd2;
		9'd347: data = 6'd0;
		9'd348: data = 6'd0;
		9'd349: data = 6'd0;
		9'd350: data = 6'd0;
		9'd351: data = 6'd0;
		9'd352: data = 6'd4;
		9'd353: data = 6'd0;
		9'd354: data = 6'd4;
		9'd355: data = 6'd0;
		9'd356: data = 6'd7;
		9'd357: data = 6'd27;
		9'd358: data = 6'd2;
		9'd359: data = 6'd0;
		9'd360: data = 6'd8;
		9'd361: data = 6'd0;
		9'd362: data = 6'd8;
		9'd363: data = 6'd0;
		9'd364: data = 6'd16;
		9'd365: data = 6'd0;
		9'd366: data = 6'd13;
		9'd367: data = 6'd6;
		9'd368: data = 6'd4;
		9'd369: data = 6'd4;
		9'd370: data = 6'd3;
		9'd371: data = 6'd3;
		9'd372: data = 6'd2;
		9'd373: data = 6'd40;
		9'd374: data = 6'd2;
		9'd375: data = 6'd0;
		9'd376: data = 6'd1;
		9'd377: data = 6'd0;
		9'd378: data = 6'd3;
		9'd379: data = 6'd2;
		9'd380: data = 6'd0;
		9'd381: data = 6'd0;
		9'd382: data = 6'd0;
		9'd383: data = 6'd0;
		9'd384: data = 6'd8;
		9'd385: data = 6'd41;
		9'd386: data = 6'd8;
		9'd387: data = 6'd0;
		9'd388: data = 6'd2;
		9'd389: data = 6'd0;
		9'd390: data = 6'd2;
		9'd391: data = 6'd0;
		9'd392: data = 6'd1;
		9'd393: data = 6'd0;
		9'd394: data = 6'd1;
		9'd395: data = 6'd0;
		9'd396: data = 6'd10;
		9'd397: data = 6'd0;
		9'd398: data = 6'd10;
		9'd399: data = 6'd0;
		9'd400: data = 6'd6;
		9'd401: data = 6'd6;
		9'd402: data = 6'd4;
		9'd403: data = 6'd6;
		9'd404: data = 6'd4;
		9'd405: data = 6'd0;
		9'd406: data = 6'd0;
		9'd407: data = 6'd0;
		9'd408: data = 6'd24;
		9'd409: data = 6'd0;
		9'd410: data = 6'd42;
		9'd411: data = 6'd0;
		9'd412: data = 6'd0;
		9'd413: data = 6'd0;
		9'd414: data = 6'd0;
		9'd415: data = 6'd0;
		9'd416: data = 6'd4;
		9'd417: data = 6'd0;
		9'd418: data = 6'd1;
		9'd419: data = 6'd0;
		9'd420: data = 6'd2;
		9'd421: data = 6'd0;
		9'd422: data = 6'd1;
		9'd423: data = 6'd0;
		9'd424: data = 6'd1;
		9'd425: data = 6'd0;
		9'd426: data = 6'd1;
		9'd427: data = 6'd0;
		9'd428: data = 6'd0;
		9'd429: data = 6'd0;
		9'd430: data = 6'd0;
		9'd431: data = 6'd0;
		9'd432: data = 6'd5;
		9'd433: data = 6'd0;
		9'd434: data = 6'd5;
		9'd435: data = 6'd0;
		9'd436: data = 6'd6;
		9'd437: data = 6'd0;
		9'd438: data = 6'd16;
		9'd439: data = 6'd0;
		9'd440: data = 6'd43;
		9'd441: data = 6'd17;
		9'd442: data = 6'd0;
		9'd443: data = 6'd0;
		9'd444: data = 6'd0;
		9'd445: data = 6'd0;
		9'd446: data = 6'd0;
		9'd447: data = 6'd0;
		9'd448: data = 6'd1;
		9'd449: data = 6'd0;
		9'd450: data = 6'd2;
		9'd451: data = 6'd0;
		9'd452: data = 6'd2;
		9'd453: data = 6'd0;
		9'd454: data = 6'd1;
		9'd455: data = 6'd0;
		9'd456: data = 6'd1;
		9'd457: data = 6'd0;
		9'd458: data = 6'd0;
		9'd459: data = 6'd0;
		9'd460: data = 6'd0;
		9'd461: data = 6'd0;
		9'd462: data = 6'd0;
		9'd463: data = 6'd0;
		9'd464: data = 6'd0;
		9'd465: data = 6'd0;
		9'd466: data = 6'd0;
		9'd467: data = 6'd0;
		9'd468: data = 6'd5;
		9'd469: data = 6'd0;
		9'd470: data = 6'd10;
		9'd471: data = 6'd17;
		9'd472: data = 6'd7;
		9'd473: data = 6'd0;
		9'd474: data = 6'd0;
		9'd475: data = 6'd1;
		9'd476: data = 6'd0;
		9'd477: data = 6'd0;
		9'd478: data = 6'd0;
		9'd479: data = 6'd0;
		9'd480: data = 6'd0;
		9'd481: data = 6'd0;
		9'd482: data = 6'd2;
		9'd483: data = 6'd0;
		9'd484: data = 6'd2;
		9'd485: data = 6'd1;
		9'd486: data = 6'd1;
		9'd487: data = 6'd1;
		9'd488: data = 6'd1;
		9'd489: data = 6'd0;
		9'd490: data = 6'd0;
		9'd491: data = 6'd0;
		9'd492: data = 6'd0;
		9'd493: data = 6'd0;
		9'd494: data = 6'd0;
		9'd495: data = 6'd0;
		9'd496: data = 6'd0;
		9'd497: data = 6'd0;
		9'd498: data = 6'd0;
		9'd499: data = 6'd0;
		9'd500: data = 6'd0;
		9'd501: data = 6'd0;
		9'd502: data = 6'd0;
		9'd503: data = 6'd0;
		9'd504: data = 6'd0;
		9'd505: data = 6'd0;
		9'd506: data = 6'd0;
		9'd507: data = 6'd2;
		9'd508: data = 6'd0;
		9'd509: data = 6'd0;
		9'd510: data = 6'd0;
		9'd511: data = 6'd0;
		default: data = 6'd0;
	endcase
end
endmodule

module layer0_N23_rsh_1(address, data);
input wire [8:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		9'd0: data = 2'd0;
		9'd1: data = 2'd0;
		9'd2: data = 2'd0;
		9'd3: data = 2'd0;
		9'd4: data = 2'd0;
		9'd5: data = 2'd0;
		9'd6: data = 2'd1;
		9'd7: data = 2'd0;
		9'd8: data = 2'd0;
		9'd9: data = 2'd0;
		9'd10: data = 2'd0;
		9'd11: data = 2'd0;
		9'd12: data = 2'd0;
		9'd13: data = 2'd0;
		9'd14: data = 2'd0;
		9'd15: data = 2'd0;
		9'd16: data = 2'd0;
		9'd17: data = 2'd0;
		9'd18: data = 2'd1;
		9'd19: data = 2'd0;
		9'd20: data = 2'd0;
		9'd21: data = 2'd0;
		9'd22: data = 2'd0;
		9'd23: data = 2'd1;
		9'd24: data = 2'd0;
		9'd25: data = 2'd1;
		9'd26: data = 2'd0;
		9'd27: data = 2'd1;
		9'd28: data = 2'd0;
		9'd29: data = 2'd1;
		9'd30: data = 2'd3;
		9'd31: data = 2'd1;
		9'd32: data = 2'd0;
		9'd33: data = 2'd0;
		9'd34: data = 2'd0;
		9'd35: data = 2'd0;
		9'd36: data = 2'd0;
		9'd37: data = 2'd3;
		9'd38: data = 2'd1;
		9'd39: data = 2'd3;
		9'd40: data = 2'd0;
		9'd41: data = 2'd1;
		9'd42: data = 2'd0;
		9'd43: data = 2'd1;
		9'd44: data = 2'd1;
		9'd45: data = 2'd1;
		9'd46: data = 2'd0;
		9'd47: data = 2'd0;
		9'd48: data = 2'd0;
		9'd49: data = 2'd0;
		9'd50: data = 2'd0;
		9'd51: data = 2'd0;
		9'd52: data = 2'd0;
		9'd53: data = 2'd1;
		9'd54: data = 2'd1;
		9'd55: data = 2'd1;
		9'd56: data = 2'd0;
		9'd57: data = 2'd1;
		9'd58: data = 2'd0;
		9'd59: data = 2'd3;
		9'd60: data = 2'd0;
		9'd61: data = 2'd0;
		9'd62: data = 2'd3;
		9'd63: data = 2'd0;
		9'd64: data = 2'd0;
		9'd65: data = 2'd3;
		9'd66: data = 2'd0;
		9'd67: data = 2'd3;
		9'd68: data = 2'd0;
		9'd69: data = 2'd3;
		9'd70: data = 2'd0;
		9'd71: data = 2'd3;
		9'd72: data = 2'd1;
		9'd73: data = 2'd1;
		9'd74: data = 2'd0;
		9'd75: data = 2'd1;
		9'd76: data = 2'd1;
		9'd77: data = 2'd0;
		9'd78: data = 2'd0;
		9'd79: data = 2'd0;
		9'd80: data = 2'd1;
		9'd81: data = 2'd0;
		9'd82: data = 2'd0;
		9'd83: data = 2'd0;
		9'd84: data = 2'd0;
		9'd85: data = 2'd0;
		9'd86: data = 2'd0;
		9'd87: data = 2'd0;
		9'd88: data = 2'd0;
		9'd89: data = 2'd3;
		9'd90: data = 2'd0;
		9'd91: data = 2'd3;
		9'd92: data = 2'd0;
		9'd93: data = 2'd3;
		9'd94: data = 2'd3;
		9'd95: data = 2'd3;
		9'd96: data = 2'd0;
		9'd97: data = 2'd3;
		9'd98: data = 2'd0;
		9'd99: data = 2'd3;
		9'd100: data = 2'd0;
		9'd101: data = 2'd3;
		9'd102: data = 2'd0;
		9'd103: data = 2'd3;
		9'd104: data = 2'd1;
		9'd105: data = 2'd1;
		9'd106: data = 2'd0;
		9'd107: data = 2'd1;
		9'd108: data = 2'd0;
		9'd109: data = 2'd1;
		9'd110: data = 2'd1;
		9'd111: data = 2'd1;
		9'd112: data = 2'd1;
		9'd113: data = 2'd1;
		9'd114: data = 2'd1;
		9'd115: data = 2'd2;
		9'd116: data = 2'd2;
		9'd117: data = 2'd3;
		9'd118: data = 2'd1;
		9'd119: data = 2'd3;
		9'd120: data = 2'd0;
		9'd121: data = 2'd3;
		9'd122: data = 2'd0;
		9'd123: data = 2'd0;
		9'd124: data = 2'd1;
		9'd125: data = 2'd1;
		9'd126: data = 2'd3;
		9'd127: data = 2'd3;
		9'd128: data = 2'd1;
		9'd129: data = 2'd3;
		9'd130: data = 2'd0;
		9'd131: data = 2'd3;
		9'd132: data = 2'd0;
		9'd133: data = 2'd3;
		9'd134: data = 2'd0;
		9'd135: data = 2'd3;
		9'd136: data = 2'd1;
		9'd137: data = 2'd1;
		9'd138: data = 2'd0;
		9'd139: data = 2'd1;
		9'd140: data = 2'd0;
		9'd141: data = 2'd1;
		9'd142: data = 2'd1;
		9'd143: data = 2'd1;
		9'd144: data = 2'd1;
		9'd145: data = 2'd1;
		9'd146: data = 2'd1;
		9'd147: data = 2'd1;
		9'd148: data = 2'd1;
		9'd149: data = 2'd1;
		9'd150: data = 2'd1;
		9'd151: data = 2'd2;
		9'd152: data = 2'd0;
		9'd153: data = 2'd0;
		9'd154: data = 2'd0;
		9'd155: data = 2'd3;
		9'd156: data = 2'd1;
		9'd157: data = 2'd0;
		9'd158: data = 2'd3;
		9'd159: data = 2'd3;
		9'd160: data = 2'd1;
		9'd161: data = 2'd3;
		9'd162: data = 2'd1;
		9'd163: data = 2'd3;
		9'd164: data = 2'd0;
		9'd165: data = 2'd3;
		9'd166: data = 2'd0;
		9'd167: data = 2'd3;
		9'd168: data = 2'd0;
		9'd169: data = 2'd1;
		9'd170: data = 2'd1;
		9'd171: data = 2'd3;
		9'd172: data = 2'd0;
		9'd173: data = 2'd3;
		9'd174: data = 2'd0;
		9'd175: data = 2'd0;
		9'd176: data = 2'd1;
		9'd177: data = 2'd1;
		9'd178: data = 2'd1;
		9'd179: data = 2'd1;
		9'd180: data = 2'd1;
		9'd181: data = 2'd1;
		9'd182: data = 2'd0;
		9'd183: data = 2'd0;
		9'd184: data = 2'd0;
		9'd185: data = 2'd3;
		9'd186: data = 2'd0;
		9'd187: data = 2'd3;
		9'd188: data = 2'd1;
		9'd189: data = 2'd3;
		9'd190: data = 2'd3;
		9'd191: data = 2'd3;
		9'd192: data = 2'd2;
		9'd193: data = 2'd3;
		9'd194: data = 2'd1;
		9'd195: data = 2'd3;
		9'd196: data = 2'd0;
		9'd197: data = 2'd3;
		9'd198: data = 2'd0;
		9'd199: data = 2'd3;
		9'd200: data = 2'd1;
		9'd201: data = 2'd2;
		9'd202: data = 2'd1;
		9'd203: data = 2'd3;
		9'd204: data = 2'd0;
		9'd205: data = 2'd3;
		9'd206: data = 2'd0;
		9'd207: data = 2'd3;
		9'd208: data = 2'd0;
		9'd209: data = 2'd0;
		9'd210: data = 2'd1;
		9'd211: data = 2'd0;
		9'd212: data = 2'd1;
		9'd213: data = 2'd3;
		9'd214: data = 2'd1;
		9'd215: data = 2'd3;
		9'd216: data = 2'd0;
		9'd217: data = 2'd3;
		9'd218: data = 2'd0;
		9'd219: data = 2'd0;
		9'd220: data = 2'd3;
		9'd221: data = 2'd2;
		9'd222: data = 2'd3;
		9'd223: data = 2'd3;
		9'd224: data = 2'd0;
		9'd225: data = 2'd0;
		9'd226: data = 2'd1;
		9'd227: data = 2'd3;
		9'd228: data = 2'd1;
		9'd229: data = 2'd3;
		9'd230: data = 2'd0;
		9'd231: data = 2'd3;
		9'd232: data = 2'd1;
		9'd233: data = 2'd1;
		9'd234: data = 2'd0;
		9'd235: data = 2'd2;
		9'd236: data = 2'd1;
		9'd237: data = 2'd2;
		9'd238: data = 2'd1;
		9'd239: data = 2'd3;
		9'd240: data = 2'd0;
		9'd241: data = 2'd3;
		9'd242: data = 2'd0;
		9'd243: data = 2'd3;
		9'd244: data = 2'd0;
		9'd245: data = 2'd3;
		9'd246: data = 2'd0;
		9'd247: data = 2'd3;
		9'd248: data = 2'd0;
		9'd249: data = 2'd0;
		9'd250: data = 2'd0;
		9'd251: data = 2'd0;
		9'd252: data = 2'd3;
		9'd253: data = 2'd1;
		9'd254: data = 2'd3;
		9'd255: data = 2'd3;
		9'd256: data = 2'd1;
		9'd257: data = 2'd0;
		9'd258: data = 2'd1;
		9'd259: data = 2'd0;
		9'd260: data = 2'd1;
		9'd261: data = 2'd3;
		9'd262: data = 2'd0;
		9'd263: data = 2'd3;
		9'd264: data = 2'd0;
		9'd265: data = 2'd0;
		9'd266: data = 2'd1;
		9'd267: data = 2'd1;
		9'd268: data = 2'd1;
		9'd269: data = 2'd1;
		9'd270: data = 2'd1;
		9'd271: data = 2'd2;
		9'd272: data = 2'd1;
		9'd273: data = 2'd2;
		9'd274: data = 2'd2;
		9'd275: data = 2'd3;
		9'd276: data = 2'd0;
		9'd277: data = 2'd3;
		9'd278: data = 2'd0;
		9'd279: data = 2'd3;
		9'd280: data = 2'd0;
		9'd281: data = 2'd0;
		9'd282: data = 2'd0;
		9'd283: data = 2'd3;
		9'd284: data = 2'd3;
		9'd285: data = 2'd0;
		9'd286: data = 2'd3;
		9'd287: data = 2'd3;
		9'd288: data = 2'd1;
		9'd289: data = 2'd3;
		9'd290: data = 2'd0;
		9'd291: data = 2'd3;
		9'd292: data = 2'd1;
		9'd293: data = 2'd3;
		9'd294: data = 2'd0;
		9'd295: data = 2'd3;
		9'd296: data = 2'd0;
		9'd297: data = 2'd3;
		9'd298: data = 2'd1;
		9'd299: data = 2'd1;
		9'd300: data = 2'd0;
		9'd301: data = 2'd1;
		9'd302: data = 2'd1;
		9'd303: data = 2'd1;
		9'd304: data = 2'd1;
		9'd305: data = 2'd1;
		9'd306: data = 2'd2;
		9'd307: data = 2'd2;
		9'd308: data = 2'd2;
		9'd309: data = 2'd2;
		9'd310: data = 2'd1;
		9'd311: data = 2'd3;
		9'd312: data = 2'd1;
		9'd313: data = 2'd0;
		9'd314: data = 2'd0;
		9'd315: data = 2'd3;
		9'd316: data = 2'd3;
		9'd317: data = 2'd3;
		9'd318: data = 2'd3;
		9'd319: data = 2'd3;
		9'd320: data = 2'd0;
		9'd321: data = 2'd0;
		9'd322: data = 2'd0;
		9'd323: data = 2'd3;
		9'd324: data = 2'd0;
		9'd325: data = 2'd3;
		9'd326: data = 2'd0;
		9'd327: data = 2'd3;
		9'd328: data = 2'd0;
		9'd329: data = 2'd3;
		9'd330: data = 2'd0;
		9'd331: data = 2'd3;
		9'd332: data = 2'd1;
		9'd333: data = 2'd1;
		9'd334: data = 2'd1;
		9'd335: data = 2'd1;
		9'd336: data = 2'd1;
		9'd337: data = 2'd1;
		9'd338: data = 2'd1;
		9'd339: data = 2'd1;
		9'd340: data = 2'd1;
		9'd341: data = 2'd1;
		9'd342: data = 2'd1;
		9'd343: data = 2'd0;
		9'd344: data = 2'd0;
		9'd345: data = 2'd3;
		9'd346: data = 2'd1;
		9'd347: data = 2'd2;
		9'd348: data = 2'd3;
		9'd349: data = 2'd3;
		9'd350: data = 2'd3;
		9'd351: data = 2'd3;
		9'd352: data = 2'd1;
		9'd353: data = 2'd3;
		9'd354: data = 2'd1;
		9'd355: data = 2'd3;
		9'd356: data = 2'd0;
		9'd357: data = 2'd0;
		9'd358: data = 2'd1;
		9'd359: data = 2'd3;
		9'd360: data = 2'd0;
		9'd361: data = 2'd3;
		9'd362: data = 2'd0;
		9'd363: data = 2'd3;
		9'd364: data = 2'd0;
		9'd365: data = 2'd3;
		9'd366: data = 2'd0;
		9'd367: data = 2'd0;
		9'd368: data = 2'd1;
		9'd369: data = 2'd1;
		9'd370: data = 2'd1;
		9'd371: data = 2'd1;
		9'd372: data = 2'd1;
		9'd373: data = 2'd0;
		9'd374: data = 2'd1;
		9'd375: data = 2'd3;
		9'd376: data = 2'd0;
		9'd377: data = 2'd3;
		9'd378: data = 2'd1;
		9'd379: data = 2'd1;
		9'd380: data = 2'd3;
		9'd381: data = 2'd3;
		9'd382: data = 2'd3;
		9'd383: data = 2'd3;
		9'd384: data = 2'd0;
		9'd385: data = 2'd0;
		9'd386: data = 2'd0;
		9'd387: data = 2'd3;
		9'd388: data = 2'd1;
		9'd389: data = 2'd3;
		9'd390: data = 2'd1;
		9'd391: data = 2'd3;
		9'd392: data = 2'd1;
		9'd393: data = 2'd3;
		9'd394: data = 2'd1;
		9'd395: data = 2'd3;
		9'd396: data = 2'd0;
		9'd397: data = 2'd3;
		9'd398: data = 2'd0;
		9'd399: data = 2'd3;
		9'd400: data = 2'd0;
		9'd401: data = 2'd0;
		9'd402: data = 2'd1;
		9'd403: data = 2'd0;
		9'd404: data = 2'd1;
		9'd405: data = 2'd3;
		9'd406: data = 2'd1;
		9'd407: data = 2'd3;
		9'd408: data = 2'd0;
		9'd409: data = 2'd3;
		9'd410: data = 2'd0;
		9'd411: data = 2'd3;
		9'd412: data = 2'd3;
		9'd413: data = 2'd3;
		9'd414: data = 2'd3;
		9'd415: data = 2'd3;
		9'd416: data = 2'd1;
		9'd417: data = 2'd3;
		9'd418: data = 2'd0;
		9'd419: data = 2'd3;
		9'd420: data = 2'd1;
		9'd421: data = 2'd2;
		9'd422: data = 2'd1;
		9'd423: data = 2'd2;
		9'd424: data = 2'd1;
		9'd425: data = 2'd3;
		9'd426: data = 2'd1;
		9'd427: data = 2'd3;
		9'd428: data = 2'd2;
		9'd429: data = 2'd3;
		9'd430: data = 2'd2;
		9'd431: data = 2'd3;
		9'd432: data = 2'd0;
		9'd433: data = 2'd3;
		9'd434: data = 2'd0;
		9'd435: data = 2'd3;
		9'd436: data = 2'd0;
		9'd437: data = 2'd3;
		9'd438: data = 2'd0;
		9'd439: data = 2'd3;
		9'd440: data = 2'd0;
		9'd441: data = 2'd0;
		9'd442: data = 2'd3;
		9'd443: data = 2'd3;
		9'd444: data = 2'd3;
		9'd445: data = 2'd3;
		9'd446: data = 2'd3;
		9'd447: data = 2'd3;
		9'd448: data = 2'd1;
		9'd449: data = 2'd3;
		9'd450: data = 2'd0;
		9'd451: data = 2'd2;
		9'd452: data = 2'd1;
		9'd453: data = 2'd2;
		9'd454: data = 2'd1;
		9'd455: data = 2'd2;
		9'd456: data = 2'd1;
		9'd457: data = 2'd2;
		9'd458: data = 2'd2;
		9'd459: data = 2'd2;
		9'd460: data = 2'd2;
		9'd461: data = 2'd3;
		9'd462: data = 2'd2;
		9'd463: data = 2'd3;
		9'd464: data = 2'd3;
		9'd465: data = 2'd3;
		9'd466: data = 2'd3;
		9'd467: data = 2'd3;
		9'd468: data = 2'd0;
		9'd469: data = 2'd3;
		9'd470: data = 2'd0;
		9'd471: data = 2'd0;
		9'd472: data = 2'd0;
		9'd473: data = 2'd3;
		9'd474: data = 2'd3;
		9'd475: data = 2'd1;
		9'd476: data = 2'd3;
		9'd477: data = 2'd3;
		9'd478: data = 2'd3;
		9'd479: data = 2'd3;
		9'd480: data = 2'd2;
		9'd481: data = 2'd3;
		9'd482: data = 2'd0;
		9'd483: data = 2'd2;
		9'd484: data = 2'd1;
		9'd485: data = 2'd1;
		9'd486: data = 2'd1;
		9'd487: data = 2'd1;
		9'd488: data = 2'd1;
		9'd489: data = 2'd2;
		9'd490: data = 2'd2;
		9'd491: data = 2'd2;
		9'd492: data = 2'd2;
		9'd493: data = 2'd2;
		9'd494: data = 2'd3;
		9'd495: data = 2'd2;
		9'd496: data = 2'd3;
		9'd497: data = 2'd3;
		9'd498: data = 2'd3;
		9'd499: data = 2'd3;
		9'd500: data = 2'd3;
		9'd501: data = 2'd3;
		9'd502: data = 2'd2;
		9'd503: data = 2'd3;
		9'd504: data = 2'd1;
		9'd505: data = 2'd3;
		9'd506: data = 2'd3;
		9'd507: data = 2'd1;
		9'd508: data = 2'd3;
		9'd509: data = 2'd3;
		9'd510: data = 2'd3;
		9'd511: data = 2'd3;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N23(address, data);
input wire [11:0] address;
output reg [3:0] data;

wire [5:0] i; layer0_N23_idx_1 idx_1_inst(address[11:3], i);
wire [1:0] t; layer0_N23_rsh_1 rsh_1_inst(address[11:3], t);
wire [3:0] b; layer0_N23_2 layer0_N23_2_inst(address[11:3], b);
wire [2:0] u; layer0_N23_ust_1 ust_1_inst({i, address[2:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule
