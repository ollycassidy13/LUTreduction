
module layer0_N6_ust_3(address, data);
input wire [5:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		6'd0: data = 2'd2;
		6'd1: data = 2'd1;
		6'd2: data = 2'd1;
		6'd3: data = 2'd0;
		6'd4: data = 2'd3;
		6'd5: data = 2'd2;
		6'd6: data = 2'd1;
		6'd7: data = 2'd1;
		6'd8: data = 2'd2;
		6'd9: data = 2'd2;
		6'd10: data = 2'd1;
		6'd11: data = 2'd1;
		6'd12: data = 2'd3;
		6'd13: data = 2'd2;
		6'd14: data = 2'd1;
		6'd15: data = 2'd1;
		6'd16: data = 2'd3;
		6'd17: data = 2'd2;
		6'd18: data = 2'd2;
		6'd19: data = 2'd1;
		6'd20: data = 2'd2;
		6'd21: data = 2'd2;
		6'd22: data = 2'd2;
		6'd23: data = 2'd1;
		6'd24: data = 2'd1;
		6'd25: data = 2'd1;
		6'd26: data = 2'd1;
		6'd27: data = 2'd1;
		6'd28: data = 2'd1;
		6'd29: data = 2'd0;
		6'd30: data = 2'd0;
		6'd31: data = 2'd1;
		6'd32: data = 2'd3;
		6'd33: data = 2'd3;
		6'd34: data = 2'd3;
		6'd35: data = 2'd3;
		6'd36: data = 2'd2;
		6'd37: data = 2'd2;
		6'd38: data = 2'd2;
		6'd39: data = 2'd2;
		6'd40: data = 2'd0;
		6'd41: data = 2'd1;
		6'd42: data = 2'd1;
		6'd43: data = 2'd2;
		6'd44: data = 2'd0;
		6'd45: data = 2'd1;
		6'd46: data = 2'd1;
		6'd47: data = 2'd2;
		6'd48: data = 2'd0;
		6'd49: data = 2'd0;
		6'd50: data = 2'd1;
		6'd51: data = 2'd2;
		6'd52: data = 2'd0;
		6'd53: data = 2'd0;
		6'd54: data = 2'd1;
		6'd55: data = 2'd1;
		6'd56: data = 2'd0;
		6'd57: data = 2'd0;
		6'd58: data = 2'd1;
		6'd59: data = 2'd1;
		6'd60: data = 2'd0;
		6'd61: data = 2'd0;
		6'd62: data = 2'd1;
		6'd63: data = 2'd1;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N6_bias_3(address, data);
input wire [0:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		1'd0: data = 2'd3;
		1'd1: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N6_idx_3(address, data);
input wire [0:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		1'd0: data = 1'd0;
		1'd1: data = 1'd1;
		default: data = 1'd0;
	endcase
end
endmodule

module layer0_N6_lb_3(address, data);
input wire [5:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		6'd0: data = 1'd0;
		6'd1: data = 1'd0;
		6'd2: data = 1'd0;
		6'd3: data = 1'd1;
		6'd4: data = 1'd0;
		6'd5: data = 1'd0;
		6'd6: data = 1'd1;
		6'd7: data = 1'd1;
		6'd8: data = 1'd1;
		6'd9: data = 1'd0;
		6'd10: data = 1'd1;
		6'd11: data = 1'd0;
		6'd12: data = 1'd0;
		6'd13: data = 1'd0;
		6'd14: data = 1'd1;
		6'd15: data = 1'd0;
		6'd16: data = 1'd0;
		6'd17: data = 1'd1;
		6'd18: data = 1'd0;
		6'd19: data = 1'd1;
		6'd20: data = 1'd1;
		6'd21: data = 1'd1;
		6'd22: data = 1'd0;
		6'd23: data = 1'd1;
		6'd24: data = 1'd1;
		6'd25: data = 1'd1;
		6'd26: data = 1'd1;
		6'd27: data = 1'd1;
		6'd28: data = 1'd0;
		6'd29: data = 1'd1;
		6'd30: data = 1'd1;
		6'd31: data = 1'd0;
		6'd32: data = 1'd1;
		6'd33: data = 1'd0;
		6'd34: data = 1'd1;
		6'd35: data = 1'd1;
		6'd36: data = 1'd0;
		6'd37: data = 1'd0;
		6'd38: data = 1'd0;
		6'd39: data = 1'd1;
		6'd40: data = 1'd1;
		6'd41: data = 1'd0;
		6'd42: data = 1'd1;
		6'd43: data = 1'd0;
		6'd44: data = 1'd0;
		6'd45: data = 1'd0;
		6'd46: data = 1'd1;
		6'd47: data = 1'd0;
		6'd48: data = 1'd0;
		6'd49: data = 1'd1;
		6'd50: data = 1'd1;
		6'd51: data = 1'd0;
		6'd52: data = 1'd0;
		6'd53: data = 1'd1;
		6'd54: data = 1'd1;
		6'd55: data = 1'd1;
		6'd56: data = 1'd0;
		6'd57: data = 1'd1;
		6'd58: data = 1'd1;
		6'd59: data = 1'd1;
		6'd60: data = 1'd0;
		6'd61: data = 1'd1;
		6'd62: data = 1'd0;
		6'd63: data = 1'd1;
		default: data = 1'd0;
	endcase
end
endmodule

module layer0_N6_3(address, data);
input wire [5:0] address;
output reg [3:0] data;

wire [0:0] i; layer0_N6_idx_3 idx_3_inst(address[5:5], i);
wire [1:0] b; layer0_N6_bias_3 bias_3_inst(address[5:5], b);
wire [0:0] lb; layer0_N6_lb_3 lb_3_inst(address, lb);
wire [1:0] u; layer0_N6_ust_3 ust_3_inst({i, address[4:0]}, u);

always @(*) begin
	data = {u + b, lb};
end
endmodule

module layer0_N6_ust_2(address, data);
input wire [7:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		8'd0: data = 2'd2;
		8'd1: data = 2'd1;
		8'd2: data = 2'd2;
		8'd3: data = 2'd1;
		8'd4: data = 2'd2;
		8'd5: data = 2'd1;
		8'd6: data = 2'd2;
		8'd7: data = 2'd0;
		8'd8: data = 2'd2;
		8'd9: data = 2'd1;
		8'd10: data = 2'd2;
		8'd11: data = 2'd1;
		8'd12: data = 2'd1;
		8'd13: data = 2'd1;
		8'd14: data = 2'd1;
		8'd15: data = 2'd0;
		8'd16: data = 2'd1;
		8'd17: data = 2'd0;
		8'd18: data = 2'd1;
		8'd19: data = 2'd1;
		8'd20: data = 2'd1;
		8'd21: data = 2'd1;
		8'd22: data = 2'd1;
		8'd23: data = 2'd1;
		8'd24: data = 2'd1;
		8'd25: data = 2'd0;
		8'd26: data = 2'd2;
		8'd27: data = 2'd1;
		8'd28: data = 2'd2;
		8'd29: data = 2'd1;
		8'd30: data = 2'd2;
		8'd31: data = 2'd1;
		8'd32: data = 2'd0;
		8'd33: data = 2'd2;
		8'd34: data = 2'd0;
		8'd35: data = 2'd2;
		8'd36: data = 2'd0;
		8'd37: data = 2'd2;
		8'd38: data = 2'd0;
		8'd39: data = 2'd2;
		8'd40: data = 2'd2;
		8'd41: data = 2'd0;
		8'd42: data = 2'd2;
		8'd43: data = 2'd0;
		8'd44: data = 2'd2;
		8'd45: data = 2'd0;
		8'd46: data = 2'd1;
		8'd47: data = 2'd0;
		8'd48: data = 2'd1;
		8'd49: data = 2'd1;
		8'd50: data = 2'd1;
		8'd51: data = 2'd1;
		8'd52: data = 2'd1;
		8'd53: data = 2'd0;
		8'd54: data = 2'd1;
		8'd55: data = 2'd0;
		8'd56: data = 2'd2;
		8'd57: data = 2'd1;
		8'd58: data = 2'd1;
		8'd59: data = 2'd1;
		8'd60: data = 2'd1;
		8'd61: data = 2'd1;
		8'd62: data = 2'd1;
		8'd63: data = 2'd0;
		8'd64: data = 2'd2;
		8'd65: data = 2'd0;
		8'd66: data = 2'd2;
		8'd67: data = 2'd0;
		8'd68: data = 2'd2;
		8'd69: data = 2'd0;
		8'd70: data = 2'd2;
		8'd71: data = 2'd0;
		8'd72: data = 2'd2;
		8'd73: data = 2'd0;
		8'd74: data = 2'd2;
		8'd75: data = 2'd1;
		8'd76: data = 2'd2;
		8'd77: data = 2'd1;
		8'd78: data = 2'd2;
		8'd79: data = 2'd1;
		8'd80: data = 2'd1;
		8'd81: data = 2'd1;
		8'd82: data = 2'd1;
		8'd83: data = 2'd1;
		8'd84: data = 2'd2;
		8'd85: data = 2'd0;
		8'd86: data = 2'd2;
		8'd87: data = 2'd0;
		8'd88: data = 2'd0;
		8'd89: data = 2'd0;
		8'd90: data = 2'd1;
		8'd91: data = 2'd0;
		8'd92: data = 2'd1;
		8'd93: data = 2'd0;
		8'd94: data = 2'd2;
		8'd95: data = 2'd1;
		8'd96: data = 2'd0;
		8'd97: data = 2'd1;
		8'd98: data = 2'd0;
		8'd99: data = 2'd1;
		8'd100: data = 2'd1;
		8'd101: data = 2'd1;
		8'd102: data = 2'd1;
		8'd103: data = 2'd1;
		8'd104: data = 2'd1;
		8'd105: data = 2'd0;
		8'd106: data = 2'd1;
		8'd107: data = 2'd0;
		8'd108: data = 2'd1;
		8'd109: data = 2'd0;
		8'd110: data = 2'd1;
		8'd111: data = 2'd1;
		8'd112: data = 2'd1;
		8'd113: data = 2'd3;
		8'd114: data = 2'd1;
		8'd115: data = 2'd3;
		8'd116: data = 2'd1;
		8'd117: data = 2'd3;
		8'd118: data = 2'd0;
		8'd119: data = 2'd2;
		8'd120: data = 2'd1;
		8'd121: data = 2'd2;
		8'd122: data = 2'd0;
		8'd123: data = 2'd2;
		8'd124: data = 2'd0;
		8'd125: data = 2'd2;
		8'd126: data = 2'd0;
		8'd127: data = 2'd2;
		8'd128: data = 2'd1;
		8'd129: data = 2'd1;
		8'd130: data = 2'd1;
		8'd131: data = 2'd1;
		8'd132: data = 2'd1;
		8'd133: data = 2'd1;
		8'd134: data = 2'd1;
		8'd135: data = 2'd0;
		8'd136: data = 2'd2;
		8'd137: data = 2'd1;
		8'd138: data = 2'd2;
		8'd139: data = 2'd0;
		8'd140: data = 2'd2;
		8'd141: data = 2'd0;
		8'd142: data = 2'd2;
		8'd143: data = 2'd0;
		8'd144: data = 2'd1;
		8'd145: data = 2'd1;
		8'd146: data = 2'd1;
		8'd147: data = 2'd1;
		8'd148: data = 2'd1;
		8'd149: data = 2'd1;
		8'd150: data = 2'd0;
		8'd151: data = 2'd0;
		8'd152: data = 2'd1;
		8'd153: data = 2'd1;
		8'd154: data = 2'd0;
		8'd155: data = 2'd0;
		8'd156: data = 2'd0;
		8'd157: data = 2'd0;
		8'd158: data = 2'd0;
		8'd159: data = 2'd0;
		8'd160: data = 2'd1;
		8'd161: data = 2'd1;
		8'd162: data = 2'd1;
		8'd163: data = 2'd0;
		8'd164: data = 2'd0;
		8'd165: data = 2'd0;
		8'd166: data = 2'd0;
		8'd167: data = 2'd0;
		8'd168: data = 2'd1;
		8'd169: data = 2'd1;
		8'd170: data = 2'd1;
		8'd171: data = 2'd0;
		8'd172: data = 2'd1;
		8'd173: data = 2'd0;
		8'd174: data = 2'd0;
		8'd175: data = 2'd0;
		8'd176: data = 2'd1;
		8'd177: data = 2'd0;
		8'd178: data = 2'd1;
		8'd179: data = 2'd0;
		8'd180: data = 2'd1;
		8'd181: data = 2'd1;
		8'd182: data = 2'd1;
		8'd183: data = 2'd0;
		8'd184: data = 2'd0;
		8'd185: data = 2'd1;
		8'd186: data = 2'd0;
		8'd187: data = 2'd1;
		8'd188: data = 2'd0;
		8'd189: data = 2'd0;
		8'd190: data = 2'd0;
		8'd191: data = 2'd0;
		8'd192: data = 2'd0;
		8'd193: data = 2'd0;
		8'd194: data = 2'd1;
		8'd195: data = 2'd0;
		8'd196: data = 2'd1;
		8'd197: data = 2'd0;
		8'd198: data = 2'd1;
		8'd199: data = 2'd1;
		8'd200: data = 2'd0;
		8'd201: data = 2'd0;
		8'd202: data = 2'd0;
		8'd203: data = 2'd0;
		8'd204: data = 2'd1;
		8'd205: data = 2'd1;
		8'd206: data = 2'd1;
		8'd207: data = 2'd1;
		8'd208: data = 2'd1;
		8'd209: data = 2'd0;
		8'd210: data = 2'd2;
		8'd211: data = 2'd0;
		8'd212: data = 2'd2;
		8'd213: data = 2'd1;
		8'd214: data = 2'd2;
		8'd215: data = 2'd1;
		8'd216: data = 2'd0;
		8'd217: data = 2'd0;
		8'd218: data = 2'd0;
		8'd219: data = 2'd0;
		8'd220: data = 2'd0;
		8'd221: data = 2'd0;
		8'd222: data = 2'd1;
		8'd223: data = 2'd1;
		8'd224: data = 2'd1;
		8'd225: data = 2'd0;
		8'd226: data = 2'd1;
		8'd227: data = 2'd0;
		8'd228: data = 2'd2;
		8'd229: data = 2'd1;
		8'd230: data = 2'd2;
		8'd231: data = 2'd1;
		8'd232: data = 2'd0;
		8'd233: data = 2'd0;
		8'd234: data = 2'd1;
		8'd235: data = 2'd0;
		8'd236: data = 2'd2;
		8'd237: data = 2'd0;
		8'd238: data = 2'd2;
		8'd239: data = 2'd1;
		8'd240: data = 2'd1;
		8'd241: data = 2'd0;
		8'd242: data = 2'd1;
		8'd243: data = 2'd1;
		8'd244: data = 2'd2;
		8'd245: data = 2'd1;
		8'd246: data = 2'd2;
		8'd247: data = 2'd1;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N6_idx_2(address, data);
input wire [5:0] address;
output reg [4:0] data;

always @(*) begin
	case(address)
		6'd0: data = 5'd4;
		6'd1: data = 5'd14;
		6'd2: data = 5'd4;
		6'd3: data = 5'd15;
		6'd4: data = 5'd1;
		6'd5: data = 5'd1;
		6'd6: data = 5'd0;
		6'd7: data = 5'd5;
		6'd8: data = 5'd16;
		6'd9: data = 5'd6;
		6'd10: data = 5'd0;
		6'd11: data = 5'd17;
		6'd12: data = 5'd0;
		6'd13: data = 5'd18;
		6'd14: data = 5'd6;
		6'd15: data = 5'd7;
		6'd16: data = 5'd0;
		6'd17: data = 5'd19;
		6'd18: data = 5'd7;
		6'd19: data = 5'd1;
		6'd20: data = 5'd0;
		6'd21: data = 5'd1;
		6'd22: data = 5'd20;
		6'd23: data = 5'd21;
		6'd24: data = 5'd8;
		6'd25: data = 5'd8;
		6'd26: data = 5'd22;
		6'd27: data = 5'd1;
		6'd28: data = 5'd5;
		6'd29: data = 5'd0;
		6'd30: data = 5'd9;
		6'd31: data = 5'd0;
		6'd32: data = 5'd0;
		6'd33: data = 5'd10;
		6'd34: data = 5'd0;
		6'd35: data = 5'd0;
		6'd36: data = 5'd0;
		6'd37: data = 5'd10;
		6'd38: data = 5'd9;
		6'd39: data = 5'd0;
		6'd40: data = 5'd23;
		6'd41: data = 5'd11;
		6'd42: data = 5'd2;
		6'd43: data = 5'd0;
		6'd44: data = 5'd12;
		6'd45: data = 5'd24;
		6'd46: data = 5'd2;
		6'd47: data = 5'd0;
		6'd48: data = 5'd12;
		6'd49: data = 5'd3;
		6'd50: data = 5'd13;
		6'd51: data = 5'd0;
		6'd52: data = 5'd25;
		6'd53: data = 5'd26;
		6'd54: data = 5'd3;
		6'd55: data = 5'd2;
		6'd56: data = 5'd27;
		6'd57: data = 5'd28;
		6'd58: data = 5'd3;
		6'd59: data = 5'd13;
		6'd60: data = 5'd11;
		6'd61: data = 5'd29;
		6'd62: data = 5'd30;
		6'd63: data = 5'd0;
		default: data = 5'd0;
	endcase
end
endmodule

module layer0_N6_rsh_2(address, data);
input wire [5:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		6'd0: data = 2'd0;
		6'd1: data = 2'd0;
		6'd2: data = 2'd0;
		6'd3: data = 2'd0;
		6'd4: data = 2'd1;
		6'd5: data = 2'd0;
		6'd6: data = 2'd0;
		6'd7: data = 2'd0;
		6'd8: data = 2'd0;
		6'd9: data = 2'd0;
		6'd10: data = 2'd1;
		6'd11: data = 2'd0;
		6'd12: data = 2'd2;
		6'd13: data = 2'd0;
		6'd14: data = 2'd0;
		6'd15: data = 2'd0;
		6'd16: data = 2'd2;
		6'd17: data = 2'd0;
		6'd18: data = 2'd1;
		6'd19: data = 2'd1;
		6'd20: data = 2'd1;
		6'd21: data = 2'd1;
		6'd22: data = 2'd0;
		6'd23: data = 2'd0;
		6'd24: data = 2'd0;
		6'd25: data = 2'd0;
		6'd26: data = 2'd0;
		6'd27: data = 2'd1;
		6'd28: data = 2'd0;
		6'd29: data = 2'd0;
		6'd30: data = 2'd0;
		6'd31: data = 2'd1;
		6'd32: data = 2'd1;
		6'd33: data = 2'd0;
		6'd34: data = 2'd1;
		6'd35: data = 2'd1;
		6'd36: data = 2'd2;
		6'd37: data = 2'd1;
		6'd38: data = 2'd0;
		6'd39: data = 2'd1;
		6'd40: data = 2'd0;
		6'd41: data = 2'd0;
		6'd42: data = 2'd0;
		6'd43: data = 2'd2;
		6'd44: data = 2'd0;
		6'd45: data = 2'd0;
		6'd46: data = 2'd0;
		6'd47: data = 2'd2;
		6'd48: data = 2'd0;
		6'd49: data = 2'd0;
		6'd50: data = 2'd0;
		6'd51: data = 2'd2;
		6'd52: data = 2'd0;
		6'd53: data = 2'd0;
		6'd54: data = 2'd1;
		6'd55: data = 2'd0;
		6'd56: data = 2'd0;
		6'd57: data = 2'd0;
		6'd58: data = 2'd1;
		6'd59: data = 2'd0;
		6'd60: data = 2'd1;
		6'd61: data = 2'd0;
		6'd62: data = 2'd0;
		6'd63: data = 2'd1;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N6_2(address, data);
input wire [8:0] address;
output reg [3:0] data;

wire [4:0] i; layer0_N6_idx_2 idx_2_inst(address[8:3], i);
wire [1:0] t; layer0_N6_rsh_2 rsh_2_inst(address[8:3], t);
wire [3:0] b; layer0_N6_3 layer0_N6_3_inst(address[8:3], b);
wire [1:0] u; layer0_N6_ust_2 ust_2_inst({i, address[2:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule

module layer0_N6_ust_1(address, data);
input wire [9:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		10'd0: data = 3'd2;
		10'd1: data = 3'd1;
		10'd2: data = 3'd1;
		10'd3: data = 3'd1;
		10'd4: data = 3'd0;
		10'd5: data = 3'd0;
		10'd6: data = 3'd0;
		10'd7: data = 3'd0;
		10'd8: data = 3'd4;
		10'd9: data = 3'd4;
		10'd10: data = 3'd3;
		10'd11: data = 3'd2;
		10'd12: data = 3'd2;
		10'd13: data = 3'd1;
		10'd14: data = 3'd0;
		10'd15: data = 3'd0;
		10'd16: data = 3'd5;
		10'd17: data = 3'd4;
		10'd18: data = 3'd4;
		10'd19: data = 3'd3;
		10'd20: data = 3'd2;
		10'd21: data = 3'd1;
		10'd22: data = 3'd0;
		10'd23: data = 3'd0;
		10'd24: data = 3'd0;
		10'd25: data = 3'd1;
		10'd26: data = 3'd1;
		10'd27: data = 3'd2;
		10'd28: data = 3'd3;
		10'd29: data = 3'd3;
		10'd30: data = 3'd4;
		10'd31: data = 3'd4;
		10'd32: data = 3'd5;
		10'd33: data = 3'd5;
		10'd34: data = 3'd5;
		10'd35: data = 3'd4;
		10'd36: data = 3'd3;
		10'd37: data = 3'd2;
		10'd38: data = 3'd1;
		10'd39: data = 3'd0;
		10'd40: data = 3'd0;
		10'd41: data = 3'd0;
		10'd42: data = 3'd0;
		10'd43: data = 3'd1;
		10'd44: data = 3'd1;
		10'd45: data = 3'd2;
		10'd46: data = 3'd3;
		10'd47: data = 3'd4;
		10'd48: data = 3'd1;
		10'd49: data = 3'd1;
		10'd50: data = 3'd1;
		10'd51: data = 3'd1;
		10'd52: data = 3'd1;
		10'd53: data = 3'd1;
		10'd54: data = 3'd1;
		10'd55: data = 3'd0;
		10'd56: data = 3'd0;
		10'd57: data = 3'd0;
		10'd58: data = 3'd1;
		10'd59: data = 3'd1;
		10'd60: data = 3'd2;
		10'd61: data = 3'd2;
		10'd62: data = 3'd3;
		10'd63: data = 3'd3;
		10'd64: data = 3'd3;
		10'd65: data = 3'd3;
		10'd66: data = 3'd3;
		10'd67: data = 3'd3;
		10'd68: data = 3'd2;
		10'd69: data = 3'd1;
		10'd70: data = 3'd0;
		10'd71: data = 3'd0;
		10'd72: data = 3'd0;
		10'd73: data = 3'd0;
		10'd74: data = 3'd0;
		10'd75: data = 3'd1;
		10'd76: data = 3'd1;
		10'd77: data = 3'd2;
		10'd78: data = 3'd2;
		10'd79: data = 3'd3;
		10'd80: data = 3'd3;
		10'd81: data = 3'd3;
		10'd82: data = 3'd3;
		10'd83: data = 3'd3;
		10'd84: data = 3'd3;
		10'd85: data = 3'd2;
		10'd86: data = 3'd1;
		10'd87: data = 3'd0;
		10'd88: data = 3'd3;
		10'd89: data = 3'd2;
		10'd90: data = 3'd1;
		10'd91: data = 3'd1;
		10'd92: data = 3'd1;
		10'd93: data = 3'd1;
		10'd94: data = 3'd0;
		10'd95: data = 3'd0;
		10'd96: data = 3'd4;
		10'd97: data = 3'd4;
		10'd98: data = 3'd4;
		10'd99: data = 3'd4;
		10'd100: data = 3'd3;
		10'd101: data = 3'd2;
		10'd102: data = 3'd1;
		10'd103: data = 3'd0;
		10'd104: data = 3'd3;
		10'd105: data = 3'd2;
		10'd106: data = 3'd2;
		10'd107: data = 3'd1;
		10'd108: data = 3'd1;
		10'd109: data = 3'd0;
		10'd110: data = 3'd0;
		10'd111: data = 3'd0;
		10'd112: data = 3'd0;
		10'd113: data = 3'd1;
		10'd114: data = 3'd2;
		10'd115: data = 3'd2;
		10'd116: data = 3'd2;
		10'd117: data = 3'd2;
		10'd118: data = 3'd2;
		10'd119: data = 3'd3;
		10'd120: data = 3'd1;
		10'd121: data = 3'd1;
		10'd122: data = 3'd1;
		10'd123: data = 3'd0;
		10'd124: data = 3'd1;
		10'd125: data = 3'd1;
		10'd126: data = 3'd1;
		10'd127: data = 3'd1;
		10'd128: data = 3'd1;
		10'd129: data = 3'd1;
		10'd130: data = 3'd0;
		10'd131: data = 3'd0;
		10'd132: data = 3'd0;
		10'd133: data = 3'd1;
		10'd134: data = 3'd1;
		10'd135: data = 3'd1;
		10'd136: data = 3'd0;
		10'd137: data = 3'd1;
		10'd138: data = 3'd1;
		10'd139: data = 3'd2;
		10'd140: data = 3'd2;
		10'd141: data = 3'd2;
		10'd142: data = 3'd2;
		10'd143: data = 3'd3;
		10'd144: data = 3'd0;
		10'd145: data = 3'd0;
		10'd146: data = 3'd1;
		10'd147: data = 3'd1;
		10'd148: data = 3'd2;
		10'd149: data = 3'd3;
		10'd150: data = 3'd4;
		10'd151: data = 3'd5;
		10'd152: data = 3'd4;
		10'd153: data = 3'd4;
		10'd154: data = 3'd3;
		10'd155: data = 3'd2;
		10'd156: data = 3'd1;
		10'd157: data = 3'd1;
		10'd158: data = 3'd0;
		10'd159: data = 3'd0;
		10'd160: data = 3'd3;
		10'd161: data = 3'd3;
		10'd162: data = 3'd2;
		10'd163: data = 3'd1;
		10'd164: data = 3'd1;
		10'd165: data = 3'd0;
		10'd166: data = 3'd0;
		10'd167: data = 3'd0;
		10'd168: data = 3'd2;
		10'd169: data = 3'd1;
		10'd170: data = 3'd1;
		10'd171: data = 3'd0;
		10'd172: data = 3'd0;
		10'd173: data = 3'd0;
		10'd174: data = 3'd0;
		10'd175: data = 3'd0;
		10'd176: data = 3'd0;
		10'd177: data = 3'd1;
		10'd178: data = 3'd1;
		10'd179: data = 3'd1;
		10'd180: data = 3'd1;
		10'd181: data = 3'd1;
		10'd182: data = 3'd1;
		10'd183: data = 3'd1;
		10'd184: data = 3'd0;
		10'd185: data = 3'd1;
		10'd186: data = 3'd1;
		10'd187: data = 3'd1;
		10'd188: data = 3'd1;
		10'd189: data = 3'd1;
		10'd190: data = 3'd1;
		10'd191: data = 3'd2;
		10'd192: data = 3'd0;
		10'd193: data = 3'd1;
		10'd194: data = 3'd2;
		10'd195: data = 3'd2;
		10'd196: data = 3'd3;
		10'd197: data = 3'd3;
		10'd198: data = 3'd3;
		10'd199: data = 3'd4;
		10'd200: data = 3'd2;
		10'd201: data = 3'd2;
		10'd202: data = 3'd2;
		10'd203: data = 3'd2;
		10'd204: data = 3'd2;
		10'd205: data = 3'd2;
		10'd206: data = 3'd1;
		10'd207: data = 3'd0;
		10'd208: data = 3'd4;
		10'd209: data = 3'd3;
		10'd210: data = 3'd3;
		10'd211: data = 3'd3;
		10'd212: data = 3'd2;
		10'd213: data = 3'd1;
		10'd214: data = 3'd0;
		10'd215: data = 3'd0;
		10'd216: data = 3'd6;
		10'd217: data = 3'd5;
		10'd218: data = 3'd5;
		10'd219: data = 3'd4;
		10'd220: data = 3'd3;
		10'd221: data = 3'd2;
		10'd222: data = 3'd1;
		10'd223: data = 3'd0;
		10'd224: data = 3'd3;
		10'd225: data = 3'd2;
		10'd226: data = 3'd2;
		10'd227: data = 3'd1;
		10'd228: data = 3'd1;
		10'd229: data = 3'd1;
		10'd230: data = 3'd0;
		10'd231: data = 3'd0;
		10'd232: data = 3'd3;
		10'd233: data = 3'd2;
		10'd234: data = 3'd2;
		10'd235: data = 3'd1;
		10'd236: data = 3'd0;
		10'd237: data = 3'd0;
		10'd238: data = 3'd0;
		10'd239: data = 3'd0;
		10'd240: data = 3'd3;
		10'd241: data = 3'd2;
		10'd242: data = 3'd1;
		10'd243: data = 3'd1;
		10'd244: data = 3'd1;
		10'd245: data = 3'd0;
		10'd246: data = 3'd0;
		10'd247: data = 3'd0;
		10'd248: data = 3'd0;
		10'd249: data = 3'd1;
		10'd250: data = 3'd1;
		10'd251: data = 3'd2;
		10'd252: data = 3'd2;
		10'd253: data = 3'd2;
		10'd254: data = 3'd3;
		10'd255: data = 3'd5;
		10'd256: data = 3'd1;
		10'd257: data = 3'd1;
		10'd258: data = 3'd1;
		10'd259: data = 3'd1;
		10'd260: data = 3'd1;
		10'd261: data = 3'd2;
		10'd262: data = 3'd1;
		10'd263: data = 3'd0;
		10'd264: data = 3'd0;
		10'd265: data = 3'd0;
		10'd266: data = 3'd0;
		10'd267: data = 3'd1;
		10'd268: data = 3'd2;
		10'd269: data = 3'd2;
		10'd270: data = 3'd2;
		10'd271: data = 3'd3;
		10'd272: data = 3'd0;
		10'd273: data = 3'd0;
		10'd274: data = 3'd0;
		10'd275: data = 3'd0;
		10'd276: data = 3'd1;
		10'd277: data = 3'd2;
		10'd278: data = 3'd3;
		10'd279: data = 3'd3;
		10'd280: data = 3'd0;
		10'd281: data = 3'd0;
		10'd282: data = 3'd1;
		10'd283: data = 3'd1;
		10'd284: data = 3'd1;
		10'd285: data = 3'd1;
		10'd286: data = 3'd1;
		10'd287: data = 3'd0;
		10'd288: data = 3'd0;
		10'd289: data = 3'd0;
		10'd290: data = 3'd1;
		10'd291: data = 3'd1;
		10'd292: data = 3'd2;
		10'd293: data = 3'd2;
		10'd294: data = 3'd2;
		10'd295: data = 3'd2;
		10'd296: data = 3'd1;
		10'd297: data = 3'd0;
		10'd298: data = 3'd0;
		10'd299: data = 3'd1;
		10'd300: data = 3'd1;
		10'd301: data = 3'd2;
		10'd302: data = 3'd3;
		10'd303: data = 3'd4;
		10'd304: data = 3'd0;
		10'd305: data = 3'd0;
		10'd306: data = 3'd1;
		10'd307: data = 3'd1;
		10'd308: data = 3'd1;
		10'd309: data = 3'd2;
		10'd310: data = 3'd2;
		10'd311: data = 3'd2;
		10'd312: data = 3'd0;
		10'd313: data = 3'd0;
		10'd314: data = 3'd0;
		10'd315: data = 3'd1;
		10'd316: data = 3'd1;
		10'd317: data = 3'd2;
		10'd318: data = 3'd3;
		10'd319: data = 3'd3;
		10'd320: data = 3'd6;
		10'd321: data = 3'd6;
		10'd322: data = 3'd5;
		10'd323: data = 3'd5;
		10'd324: data = 3'd4;
		10'd325: data = 3'd3;
		10'd326: data = 3'd2;
		10'd327: data = 3'd0;
		10'd328: data = 3'd4;
		10'd329: data = 3'd4;
		10'd330: data = 3'd4;
		10'd331: data = 3'd3;
		10'd332: data = 3'd3;
		10'd333: data = 3'd2;
		10'd334: data = 3'd1;
		10'd335: data = 3'd0;
		10'd336: data = 3'd3;
		10'd337: data = 3'd3;
		10'd338: data = 3'd2;
		10'd339: data = 3'd2;
		10'd340: data = 3'd1;
		10'd341: data = 3'd0;
		10'd342: data = 3'd0;
		10'd343: data = 3'd0;
		10'd344: data = 3'd3;
		10'd345: data = 3'd2;
		10'd346: data = 3'd2;
		10'd347: data = 3'd2;
		10'd348: data = 3'd1;
		10'd349: data = 3'd0;
		10'd350: data = 3'd0;
		10'd351: data = 3'd0;
		10'd352: data = 3'd2;
		10'd353: data = 3'd2;
		10'd354: data = 3'd2;
		10'd355: data = 3'd2;
		10'd356: data = 3'd1;
		10'd357: data = 3'd0;
		10'd358: data = 3'd0;
		10'd359: data = 3'd0;
		10'd360: data = 3'd2;
		10'd361: data = 3'd2;
		10'd362: data = 3'd2;
		10'd363: data = 3'd1;
		10'd364: data = 3'd1;
		10'd365: data = 3'd1;
		10'd366: data = 3'd1;
		10'd367: data = 3'd0;
		10'd368: data = 3'd2;
		10'd369: data = 3'd1;
		10'd370: data = 3'd1;
		10'd371: data = 3'd1;
		10'd372: data = 3'd1;
		10'd373: data = 3'd1;
		10'd374: data = 3'd1;
		10'd375: data = 3'd0;
		10'd376: data = 3'd2;
		10'd377: data = 3'd1;
		10'd378: data = 3'd1;
		10'd379: data = 3'd1;
		10'd380: data = 3'd1;
		10'd381: data = 3'd1;
		10'd382: data = 3'd0;
		10'd383: data = 3'd0;
		10'd384: data = 3'd2;
		10'd385: data = 3'd2;
		10'd386: data = 3'd1;
		10'd387: data = 3'd1;
		10'd388: data = 3'd1;
		10'd389: data = 3'd1;
		10'd390: data = 3'd0;
		10'd391: data = 3'd0;
		10'd392: data = 3'd1;
		10'd393: data = 3'd0;
		10'd394: data = 3'd0;
		10'd395: data = 3'd0;
		10'd396: data = 3'd0;
		10'd397: data = 3'd0;
		10'd398: data = 3'd0;
		10'd399: data = 3'd1;
		10'd400: data = 3'd1;
		10'd401: data = 3'd0;
		10'd402: data = 3'd0;
		10'd403: data = 3'd0;
		10'd404: data = 3'd0;
		10'd405: data = 3'd1;
		10'd406: data = 3'd1;
		10'd407: data = 3'd1;
		10'd408: data = 3'd0;
		10'd409: data = 3'd0;
		10'd410: data = 3'd1;
		10'd411: data = 3'd2;
		10'd412: data = 3'd2;
		10'd413: data = 3'd3;
		10'd414: data = 3'd4;
		10'd415: data = 3'd4;
		10'd416: data = 3'd0;
		10'd417: data = 3'd1;
		10'd418: data = 3'd2;
		10'd419: data = 3'd2;
		10'd420: data = 3'd3;
		10'd421: data = 3'd3;
		10'd422: data = 3'd4;
		10'd423: data = 3'd5;
		10'd424: data = 3'd0;
		10'd425: data = 3'd1;
		10'd426: data = 3'd1;
		10'd427: data = 3'd2;
		10'd428: data = 3'd2;
		10'd429: data = 3'd3;
		10'd430: data = 3'd4;
		10'd431: data = 3'd5;
		10'd432: data = 3'd0;
		10'd433: data = 3'd0;
		10'd434: data = 3'd1;
		10'd435: data = 3'd1;
		10'd436: data = 3'd2;
		10'd437: data = 3'd2;
		10'd438: data = 3'd3;
		10'd439: data = 3'd5;
		10'd440: data = 3'd1;
		10'd441: data = 3'd0;
		10'd442: data = 3'd0;
		10'd443: data = 3'd0;
		10'd444: data = 3'd1;
		10'd445: data = 3'd1;
		10'd446: data = 3'd1;
		10'd447: data = 3'd2;
		10'd448: data = 3'd0;
		10'd449: data = 3'd1;
		10'd450: data = 3'd1;
		10'd451: data = 3'd1;
		10'd452: data = 3'd2;
		10'd453: data = 3'd2;
		10'd454: data = 3'd3;
		10'd455: data = 3'd4;
		10'd456: data = 3'd0;
		10'd457: data = 3'd1;
		10'd458: data = 3'd1;
		10'd459: data = 3'd1;
		10'd460: data = 3'd2;
		10'd461: data = 3'd2;
		10'd462: data = 3'd2;
		10'd463: data = 3'd4;
		10'd464: data = 3'd0;
		10'd465: data = 3'd0;
		10'd466: data = 3'd1;
		10'd467: data = 3'd1;
		10'd468: data = 3'd1;
		10'd469: data = 3'd1;
		10'd470: data = 3'd1;
		10'd471: data = 3'd3;
		10'd472: data = 3'd1;
		10'd473: data = 3'd0;
		10'd474: data = 3'd1;
		10'd475: data = 3'd1;
		10'd476: data = 3'd2;
		10'd477: data = 3'd2;
		10'd478: data = 3'd3;
		10'd479: data = 3'd4;
		10'd480: data = 3'd0;
		10'd481: data = 3'd0;
		10'd482: data = 3'd0;
		10'd483: data = 3'd0;
		10'd484: data = 3'd1;
		10'd485: data = 3'd1;
		10'd486: data = 3'd3;
		10'd487: data = 3'd3;
		10'd488: data = 3'd1;
		10'd489: data = 3'd0;
		10'd490: data = 3'd1;
		10'd491: data = 3'd1;
		10'd492: data = 3'd1;
		10'd493: data = 3'd2;
		10'd494: data = 3'd3;
		10'd495: data = 3'd4;
		10'd496: data = 3'd1;
		10'd497: data = 3'd0;
		10'd498: data = 3'd0;
		10'd499: data = 3'd1;
		10'd500: data = 3'd1;
		10'd501: data = 3'd1;
		10'd502: data = 3'd3;
		10'd503: data = 3'd4;
		10'd504: data = 3'd1;
		10'd505: data = 3'd0;
		10'd506: data = 3'd0;
		10'd507: data = 3'd1;
		10'd508: data = 3'd1;
		10'd509: data = 3'd1;
		10'd510: data = 3'd2;
		10'd511: data = 3'd4;
		10'd512: data = 3'd1;
		10'd513: data = 3'd0;
		10'd514: data = 3'd0;
		10'd515: data = 3'd0;
		10'd516: data = 3'd1;
		10'd517: data = 3'd1;
		10'd518: data = 3'd2;
		10'd519: data = 3'd4;
		10'd520: data = 3'd1;
		10'd521: data = 3'd0;
		10'd522: data = 3'd0;
		10'd523: data = 3'd0;
		10'd524: data = 3'd0;
		10'd525: data = 3'd1;
		10'd526: data = 3'd1;
		10'd527: data = 3'd3;
		10'd528: data = 3'd0;
		10'd529: data = 3'd0;
		10'd530: data = 3'd0;
		10'd531: data = 3'd0;
		10'd532: data = 3'd1;
		10'd533: data = 3'd1;
		10'd534: data = 3'd2;
		10'd535: data = 3'd1;
		10'd536: data = 3'd0;
		10'd537: data = 3'd1;
		10'd538: data = 3'd1;
		10'd539: data = 3'd1;
		10'd540: data = 3'd2;
		10'd541: data = 3'd2;
		10'd542: data = 3'd2;
		10'd543: data = 3'd2;
		10'd544: data = 3'd0;
		10'd545: data = 3'd0;
		10'd546: data = 3'd0;
		10'd547: data = 3'd1;
		10'd548: data = 3'd2;
		10'd549: data = 3'd2;
		10'd550: data = 3'd2;
		10'd551: data = 3'd2;
		10'd552: data = 3'd0;
		10'd553: data = 3'd0;
		10'd554: data = 3'd1;
		10'd555: data = 3'd2;
		10'd556: data = 3'd2;
		10'd557: data = 3'd3;
		10'd558: data = 3'd3;
		10'd559: data = 3'd3;
		10'd560: data = 3'd0;
		10'd561: data = 3'd0;
		10'd562: data = 3'd0;
		10'd563: data = 3'd1;
		10'd564: data = 3'd2;
		10'd565: data = 3'd3;
		10'd566: data = 3'd3;
		10'd567: data = 3'd3;
		10'd568: data = 3'd5;
		10'd569: data = 3'd5;
		10'd570: data = 3'd5;
		10'd571: data = 3'd5;
		10'd572: data = 3'd3;
		10'd573: data = 3'd2;
		10'd574: data = 3'd1;
		10'd575: data = 3'd0;
		10'd576: data = 3'd0;
		10'd577: data = 3'd0;
		10'd578: data = 3'd1;
		10'd579: data = 3'd1;
		10'd580: data = 3'd2;
		10'd581: data = 3'd3;
		10'd582: data = 3'd4;
		10'd583: data = 3'd4;
		10'd584: data = 3'd0;
		10'd585: data = 3'd0;
		10'd586: data = 3'd1;
		10'd587: data = 3'd1;
		10'd588: data = 3'd2;
		10'd589: data = 3'd3;
		10'd590: data = 3'd3;
		10'd591: data = 3'd4;
		10'd592: data = 3'd0;
		10'd593: data = 3'd0;
		10'd594: data = 3'd0;
		10'd595: data = 3'd1;
		10'd596: data = 3'd1;
		10'd597: data = 3'd3;
		10'd598: data = 3'd3;
		10'd599: data = 3'd4;
		10'd600: data = 3'd1;
		10'd601: data = 3'd0;
		10'd602: data = 3'd1;
		10'd603: data = 3'd1;
		10'd604: data = 3'd2;
		10'd605: data = 3'd2;
		10'd606: data = 3'd4;
		10'd607: data = 3'd4;
		10'd608: data = 3'd4;
		10'd609: data = 3'd4;
		10'd610: data = 3'd5;
		10'd611: data = 3'd4;
		10'd612: data = 3'd3;
		10'd613: data = 3'd2;
		10'd614: data = 3'd1;
		10'd615: data = 3'd0;
		10'd616: data = 3'd3;
		10'd617: data = 3'd4;
		10'd618: data = 3'd4;
		10'd619: data = 3'd4;
		10'd620: data = 3'd3;
		10'd621: data = 3'd2;
		10'd622: data = 3'd1;
		10'd623: data = 3'd0;
		10'd624: data = 3'd3;
		10'd625: data = 3'd3;
		10'd626: data = 3'd3;
		10'd627: data = 3'd3;
		10'd628: data = 3'd2;
		10'd629: data = 3'd1;
		10'd630: data = 3'd1;
		10'd631: data = 3'd0;
		10'd632: data = 3'd0;
		10'd633: data = 3'd1;
		10'd634: data = 3'd1;
		10'd635: data = 3'd1;
		10'd636: data = 3'd1;
		10'd637: data = 3'd2;
		10'd638: data = 3'd2;
		10'd639: data = 3'd2;
		10'd640: data = 3'd4;
		10'd641: data = 3'd4;
		10'd642: data = 3'd4;
		10'd643: data = 3'd3;
		10'd644: data = 3'd2;
		10'd645: data = 3'd1;
		10'd646: data = 3'd0;
		10'd647: data = 3'd0;
		10'd648: data = 3'd1;
		10'd649: data = 3'd0;
		10'd650: data = 3'd1;
		10'd651: data = 3'd1;
		10'd652: data = 3'd2;
		10'd653: data = 3'd3;
		10'd654: data = 3'd3;
		10'd655: data = 3'd4;
		10'd656: data = 3'd0;
		10'd657: data = 3'd0;
		10'd658: data = 3'd1;
		10'd659: data = 3'd1;
		10'd660: data = 3'd2;
		10'd661: data = 3'd3;
		10'd662: data = 3'd3;
		10'd663: data = 3'd3;
		10'd664: data = 3'd6;
		10'd665: data = 3'd6;
		10'd666: data = 3'd5;
		10'd667: data = 3'd5;
		10'd668: data = 3'd3;
		10'd669: data = 3'd2;
		10'd670: data = 3'd1;
		10'd671: data = 3'd0;
		10'd672: data = 3'd0;
		10'd673: data = 3'd0;
		10'd674: data = 3'd0;
		10'd675: data = 3'd0;
		10'd676: data = 3'd1;
		10'd677: data = 3'd2;
		10'd678: data = 3'd2;
		10'd679: data = 3'd3;
		10'd680: data = 3'd6;
		10'd681: data = 3'd6;
		10'd682: data = 3'd5;
		10'd683: data = 3'd4;
		10'd684: data = 3'd3;
		10'd685: data = 3'd2;
		10'd686: data = 3'd1;
		10'd687: data = 3'd0;
		10'd688: data = 3'd1;
		10'd689: data = 3'd0;
		10'd690: data = 3'd0;
		10'd691: data = 3'd1;
		10'd692: data = 3'd2;
		10'd693: data = 3'd2;
		10'd694: data = 3'd3;
		10'd695: data = 3'd4;
		10'd696: data = 3'd3;
		10'd697: data = 3'd3;
		10'd698: data = 3'd3;
		10'd699: data = 3'd2;
		10'd700: data = 3'd1;
		10'd701: data = 3'd0;
		10'd702: data = 3'd0;
		10'd703: data = 3'd0;
		10'd704: data = 3'd3;
		10'd705: data = 3'd3;
		10'd706: data = 3'd3;
		10'd707: data = 3'd2;
		10'd708: data = 3'd2;
		10'd709: data = 3'd1;
		10'd710: data = 3'd0;
		10'd711: data = 3'd0;
		10'd712: data = 3'd4;
		10'd713: data = 3'd4;
		10'd714: data = 3'd4;
		10'd715: data = 3'd3;
		10'd716: data = 3'd2;
		10'd717: data = 3'd1;
		10'd718: data = 3'd1;
		10'd719: data = 3'd0;
		10'd720: data = 3'd5;
		10'd721: data = 3'd4;
		10'd722: data = 3'd4;
		10'd723: data = 3'd3;
		10'd724: data = 3'd2;
		10'd725: data = 3'd2;
		10'd726: data = 3'd0;
		10'd727: data = 3'd0;
		10'd728: data = 3'd1;
		10'd729: data = 3'd0;
		10'd730: data = 3'd1;
		10'd731: data = 3'd1;
		10'd732: data = 3'd2;
		10'd733: data = 3'd2;
		10'd734: data = 3'd3;
		10'd735: data = 3'd3;
		10'd736: data = 3'd5;
		10'd737: data = 3'd5;
		10'd738: data = 3'd4;
		10'd739: data = 3'd3;
		10'd740: data = 3'd2;
		10'd741: data = 3'd1;
		10'd742: data = 3'd0;
		10'd743: data = 3'd0;
		10'd744: data = 3'd0;
		10'd745: data = 3'd0;
		10'd746: data = 3'd0;
		10'd747: data = 3'd1;
		10'd748: data = 3'd1;
		10'd749: data = 3'd2;
		10'd750: data = 3'd2;
		10'd751: data = 3'd2;
		10'd752: data = 3'd1;
		10'd753: data = 3'd1;
		10'd754: data = 3'd1;
		10'd755: data = 3'd0;
		10'd756: data = 3'd1;
		10'd757: data = 3'd0;
		10'd758: data = 3'd0;
		10'd759: data = 3'd0;
		10'd760: data = 3'd4;
		10'd761: data = 3'd4;
		10'd762: data = 3'd3;
		10'd763: data = 3'd2;
		10'd764: data = 3'd1;
		10'd765: data = 3'd0;
		10'd766: data = 3'd0;
		10'd767: data = 3'd0;
		10'd768: data = 3'd1;
		10'd769: data = 3'd0;
		10'd770: data = 3'd0;
		10'd771: data = 3'd1;
		10'd772: data = 3'd1;
		10'd773: data = 3'd1;
		10'd774: data = 3'd1;
		10'd775: data = 3'd2;
		10'd776: data = 3'd5;
		10'd777: data = 3'd4;
		10'd778: data = 3'd3;
		10'd779: data = 3'd2;
		10'd780: data = 3'd1;
		10'd781: data = 3'd0;
		10'd782: data = 3'd0;
		10'd783: data = 3'd0;
		10'd784: data = 3'd5;
		10'd785: data = 3'd5;
		10'd786: data = 3'd4;
		10'd787: data = 3'd3;
		10'd788: data = 3'd2;
		10'd789: data = 3'd1;
		10'd790: data = 3'd1;
		10'd791: data = 3'd0;
		10'd792: data = 3'd2;
		10'd793: data = 3'd2;
		10'd794: data = 3'd1;
		10'd795: data = 3'd1;
		10'd796: data = 3'd1;
		10'd797: data = 3'd1;
		10'd798: data = 3'd1;
		10'd799: data = 3'd0;
		10'd800: data = 3'd1;
		10'd801: data = 3'd1;
		10'd802: data = 3'd0;
		10'd803: data = 3'd0;
		10'd804: data = 3'd0;
		10'd805: data = 3'd0;
		10'd806: data = 3'd0;
		10'd807: data = 3'd1;
		10'd808: data = 3'd4;
		10'd809: data = 3'd4;
		10'd810: data = 3'd3;
		10'd811: data = 3'd2;
		10'd812: data = 3'd1;
		10'd813: data = 3'd1;
		10'd814: data = 3'd1;
		10'd815: data = 3'd0;
		10'd816: data = 3'd2;
		10'd817: data = 3'd1;
		10'd818: data = 3'd2;
		10'd819: data = 3'd2;
		10'd820: data = 3'd1;
		10'd821: data = 3'd1;
		10'd822: data = 3'd1;
		10'd823: data = 3'd0;
		10'd824: data = 3'd1;
		10'd825: data = 3'd0;
		10'd826: data = 3'd0;
		10'd827: data = 3'd1;
		10'd828: data = 3'd0;
		10'd829: data = 3'd0;
		10'd830: data = 3'd0;
		10'd831: data = 3'd0;
		10'd832: data = 3'd1;
		10'd833: data = 3'd1;
		10'd834: data = 3'd1;
		10'd835: data = 3'd1;
		10'd836: data = 3'd0;
		10'd837: data = 3'd0;
		10'd838: data = 3'd1;
		10'd839: data = 3'd1;
		10'd840: data = 3'd1;
		10'd841: data = 3'd1;
		10'd842: data = 3'd1;
		10'd843: data = 3'd1;
		10'd844: data = 3'd0;
		10'd845: data = 3'd1;
		10'd846: data = 3'd1;
		10'd847: data = 3'd0;
		10'd848: data = 3'd1;
		10'd849: data = 3'd0;
		10'd850: data = 3'd1;
		10'd851: data = 3'd0;
		10'd852: data = 3'd0;
		10'd853: data = 3'd0;
		10'd854: data = 3'd0;
		10'd855: data = 3'd0;
		10'd856: data = 3'd3;
		10'd857: data = 3'd2;
		10'd858: data = 3'd2;
		10'd859: data = 3'd2;
		10'd860: data = 3'd1;
		10'd861: data = 3'd1;
		10'd862: data = 3'd1;
		10'd863: data = 3'd0;
		10'd864: data = 3'd2;
		10'd865: data = 3'd1;
		10'd866: data = 3'd1;
		10'd867: data = 3'd0;
		10'd868: data = 3'd0;
		10'd869: data = 3'd1;
		10'd870: data = 3'd1;
		10'd871: data = 3'd1;
		10'd872: data = 3'd0;
		10'd873: data = 3'd0;
		10'd874: data = 3'd0;
		10'd875: data = 3'd0;
		10'd876: data = 3'd1;
		10'd877: data = 3'd1;
		10'd878: data = 3'd1;
		10'd879: data = 3'd0;
		10'd880: data = 3'd1;
		10'd881: data = 3'd1;
		10'd882: data = 3'd0;
		10'd883: data = 3'd0;
		10'd884: data = 3'd1;
		10'd885: data = 3'd0;
		10'd886: data = 3'd0;
		10'd887: data = 3'd0;
		10'd888: data = 3'd1;
		10'd889: data = 3'd1;
		10'd890: data = 3'd0;
		10'd891: data = 3'd0;
		10'd892: data = 3'd1;
		10'd893: data = 3'd1;
		10'd894: data = 3'd1;
		10'd895: data = 3'd1;
		10'd896: data = 3'd1;
		10'd897: data = 3'd0;
		10'd898: data = 3'd0;
		10'd899: data = 3'd0;
		10'd900: data = 3'd0;
		10'd901: data = 3'd0;
		10'd902: data = 3'd1;
		10'd903: data = 3'd1;
		default: data = 3'd0;
	endcase
end
endmodule

module layer0_N6_idx_1(address, data);
input wire [8:0] address;
output reg [6:0] data;

always @(*) begin
	case(address)
		9'd0: data = 7'd23;
		9'd1: data = 7'd14;
		9'd2: data = 7'd31;
		9'd3: data = 7'd14;
		9'd4: data = 7'd3;
		9'd5: data = 7'd14;
		9'd6: data = 7'd5;
		9'd7: data = 7'd17;
		9'd8: data = 7'd24;
		9'd9: data = 7'd24;
		9'd10: data = 7'd3;
		9'd11: data = 7'd3;
		9'd12: data = 7'd3;
		9'd13: data = 7'd51;
		9'd14: data = 7'd23;
		9'd15: data = 7'd52;
		9'd16: data = 7'd5;
		9'd17: data = 7'd53;
		9'd18: data = 7'd3;
		9'd19: data = 7'd18;
		9'd20: data = 7'd3;
		9'd21: data = 7'd54;
		9'd22: data = 7'd3;
		9'd23: data = 7'd5;
		9'd24: data = 7'd5;
		9'd25: data = 7'd31;
		9'd26: data = 7'd55;
		9'd27: data = 7'd56;
		9'd28: data = 7'd5;
		9'd29: data = 7'd57;
		9'd30: data = 7'd3;
		9'd31: data = 7'd58;
		9'd32: data = 7'd32;
		9'd33: data = 7'd3;
		9'd34: data = 7'd6;
		9'd35: data = 7'd3;
		9'd36: data = 7'd25;
		9'd37: data = 7'd3;
		9'd38: data = 7'd25;
		9'd39: data = 7'd3;
		9'd40: data = 7'd6;
		9'd41: data = 7'd7;
		9'd42: data = 7'd6;
		9'd43: data = 7'd33;
		9'd44: data = 7'd25;
		9'd45: data = 7'd9;
		9'd46: data = 7'd32;
		9'd47: data = 7'd59;
		9'd48: data = 7'd6;
		9'd49: data = 7'd5;
		9'd50: data = 7'd6;
		9'd51: data = 7'd34;
		9'd52: data = 7'd6;
		9'd53: data = 7'd60;
		9'd54: data = 7'd6;
		9'd55: data = 7'd61;
		9'd56: data = 7'd6;
		9'd57: data = 7'd62;
		9'd58: data = 7'd0;
		9'd59: data = 7'd63;
		9'd60: data = 7'd0;
		9'd61: data = 7'd64;
		9'd62: data = 7'd35;
		9'd63: data = 7'd65;
		9'd64: data = 7'd10;
		9'd65: data = 7'd3;
		9'd66: data = 7'd10;
		9'd67: data = 7'd18;
		9'd68: data = 7'd10;
		9'd69: data = 7'd66;
		9'd70: data = 7'd10;
		9'd71: data = 7'd67;
		9'd72: data = 7'd12;
		9'd73: data = 7'd36;
		9'd74: data = 7'd12;
		9'd75: data = 7'd68;
		9'd76: data = 7'd12;
		9'd77: data = 7'd69;
		9'd78: data = 7'd12;
		9'd79: data = 7'd70;
		9'd80: data = 7'd71;
		9'd81: data = 7'd72;
		9'd82: data = 7'd4;
		9'd83: data = 7'd73;
		9'd84: data = 7'd4;
		9'd85: data = 7'd74;
		9'd86: data = 7'd4;
		9'd87: data = 7'd5;
		9'd88: data = 7'd4;
		9'd89: data = 7'd34;
		9'd90: data = 7'd4;
		9'd91: data = 7'd75;
		9'd92: data = 7'd76;
		9'd93: data = 7'd37;
		9'd94: data = 7'd77;
		9'd95: data = 7'd37;
		9'd96: data = 7'd8;
		9'd97: data = 7'd7;
		9'd98: data = 7'd8;
		9'd99: data = 7'd7;
		9'd100: data = 7'd78;
		9'd101: data = 7'd7;
		9'd102: data = 7'd8;
		9'd103: data = 7'd7;
		9'd104: data = 7'd12;
		9'd105: data = 7'd79;
		9'd106: data = 7'd12;
		9'd107: data = 7'd38;
		9'd108: data = 7'd80;
		9'd109: data = 7'd3;
		9'd110: data = 7'd4;
		9'd111: data = 7'd7;
		9'd112: data = 7'd4;
		9'd113: data = 7'd33;
		9'd114: data = 7'd4;
		9'd115: data = 7'd9;
		9'd116: data = 7'd4;
		9'd117: data = 7'd81;
		9'd118: data = 7'd4;
		9'd119: data = 7'd82;
		9'd120: data = 7'd4;
		9'd121: data = 7'd39;
		9'd122: data = 7'd40;
		9'd123: data = 7'd39;
		9'd124: data = 7'd83;
		9'd125: data = 7'd84;
		9'd126: data = 7'd85;
		9'd127: data = 7'd86;
		9'd128: data = 7'd87;
		9'd129: data = 7'd7;
		9'd130: data = 7'd8;
		9'd131: data = 7'd7;
		9'd132: data = 7'd8;
		9'd133: data = 7'd9;
		9'd134: data = 7'd8;
		9'd135: data = 7'd9;
		9'd136: data = 7'd88;
		9'd137: data = 7'd3;
		9'd138: data = 7'd89;
		9'd139: data = 7'd23;
		9'd140: data = 7'd26;
		9'd141: data = 7'd24;
		9'd142: data = 7'd26;
		9'd143: data = 7'd17;
		9'd144: data = 7'd8;
		9'd145: data = 7'd36;
		9'd146: data = 7'd41;
		9'd147: data = 7'd38;
		9'd148: data = 7'd90;
		9'd149: data = 7'd9;
		9'd150: data = 7'd2;
		9'd151: data = 7'd18;
		9'd152: data = 7'd2;
		9'd153: data = 7'd91;
		9'd154: data = 7'd92;
		9'd155: data = 7'd9;
		9'd156: data = 7'd27;
		9'd157: data = 7'd93;
		9'd158: data = 7'd27;
		9'd159: data = 7'd18;
		9'd160: data = 7'd42;
		9'd161: data = 7'd94;
		9'd162: data = 7'd42;
		9'd163: data = 7'd8;
		9'd164: data = 7'd43;
		9'd165: data = 7'd8;
		9'd166: data = 7'd44;
		9'd167: data = 7'd4;
		9'd168: data = 7'd2;
		9'd169: data = 7'd4;
		9'd170: data = 7'd19;
		9'd171: data = 7'd4;
		9'd172: data = 7'd43;
		9'd173: data = 7'd0;
		9'd174: data = 7'd44;
		9'd175: data = 7'd0;
		9'd176: data = 7'd13;
		9'd177: data = 7'd0;
		9'd178: data = 7'd13;
		9'd179: data = 7'd14;
		9'd180: data = 7'd1;
		9'd181: data = 7'd17;
		9'd182: data = 7'd19;
		9'd183: data = 7'd7;
		9'd184: data = 7'd19;
		9'd185: data = 7'd3;
		9'd186: data = 7'd95;
		9'd187: data = 7'd96;
		9'd188: data = 7'd97;
		9'd189: data = 7'd17;
		9'd190: data = 7'd98;
		9'd191: data = 7'd7;
		9'd192: data = 7'd45;
		9'd193: data = 7'd2;
		9'd194: data = 7'd99;
		9'd195: data = 7'd2;
		9'd196: data = 7'd46;
		9'd197: data = 7'd2;
		9'd198: data = 7'd47;
		9'd199: data = 7'd2;
		9'd200: data = 7'd10;
		9'd201: data = 7'd2;
		9'd202: data = 7'd4;
		9'd203: data = 7'd1;
		9'd204: data = 7'd2;
		9'd205: data = 7'd1;
		9'd206: data = 7'd2;
		9'd207: data = 7'd26;
		9'd208: data = 7'd28;
		9'd209: data = 7'd10;
		9'd210: data = 7'd13;
		9'd211: data = 7'd6;
		9'd212: data = 7'd20;
		9'd213: data = 7'd0;
		9'd214: data = 7'd20;
		9'd215: data = 7'd100;
		9'd216: data = 7'd20;
		9'd217: data = 7'd0;
		9'd218: data = 7'd20;
		9'd219: data = 7'd0;
		9'd220: data = 7'd101;
		9'd221: data = 7'd0;
		9'd222: data = 7'd19;
		9'd223: data = 7'd0;
		9'd224: data = 7'd1;
		9'd225: data = 7'd21;
		9'd226: data = 7'd1;
		9'd227: data = 7'd21;
		9'd228: data = 7'd0;
		9'd229: data = 7'd2;
		9'd230: data = 7'd6;
		9'd231: data = 7'd2;
		9'd232: data = 7'd10;
		9'd233: data = 7'd2;
		9'd234: data = 7'd1;
		9'd235: data = 7'd2;
		9'd236: data = 7'd1;
		9'd237: data = 7'd1;
		9'd238: data = 7'd1;
		9'd239: data = 7'd4;
		9'd240: data = 7'd2;
		9'd241: data = 7'd102;
		9'd242: data = 7'd28;
		9'd243: data = 7'd103;
		9'd244: data = 7'd28;
		9'd245: data = 7'd1;
		9'd246: data = 7'd13;
		9'd247: data = 7'd2;
		9'd248: data = 7'd13;
		9'd249: data = 7'd1;
		9'd250: data = 7'd29;
		9'd251: data = 7'd1;
		9'd252: data = 7'd29;
		9'd253: data = 7'd1;
		9'd254: data = 7'd29;
		9'd255: data = 7'd0;
		9'd256: data = 7'd1;
		9'd257: data = 7'd0;
		9'd258: data = 7'd0;
		9'd259: data = 7'd0;
		9'd260: data = 7'd0;
		9'd261: data = 7'd0;
		9'd262: data = 7'd0;
		9'd263: data = 7'd0;
		9'd264: data = 7'd48;
		9'd265: data = 7'd0;
		9'd266: data = 7'd27;
		9'd267: data = 7'd0;
		9'd268: data = 7'd0;
		9'd269: data = 7'd104;
		9'd270: data = 7'd1;
		9'd271: data = 7'd105;
		9'd272: data = 7'd1;
		9'd273: data = 7'd106;
		9'd274: data = 7'd41;
		9'd275: data = 7'd0;
		9'd276: data = 7'd11;
		9'd277: data = 7'd1;
		9'd278: data = 7'd11;
		9'd279: data = 7'd1;
		9'd280: data = 7'd11;
		9'd281: data = 7'd1;
		9'd282: data = 7'd30;
		9'd283: data = 7'd1;
		9'd284: data = 7'd30;
		9'd285: data = 7'd1;
		9'd286: data = 7'd30;
		9'd287: data = 7'd0;
		9'd288: data = 7'd2;
		9'd289: data = 7'd0;
		9'd290: data = 7'd1;
		9'd291: data = 7'd0;
		9'd292: data = 7'd2;
		9'd293: data = 7'd0;
		9'd294: data = 7'd0;
		9'd295: data = 7'd0;
		9'd296: data = 7'd13;
		9'd297: data = 7'd0;
		9'd298: data = 7'd40;
		9'd299: data = 7'd0;
		9'd300: data = 7'd45;
		9'd301: data = 7'd0;
		9'd302: data = 7'd107;
		9'd303: data = 7'd2;
		9'd304: data = 7'd0;
		9'd305: data = 7'd4;
		9'd306: data = 7'd1;
		9'd307: data = 7'd0;
		9'd308: data = 7'd48;
		9'd309: data = 7'd0;
		9'd310: data = 7'd11;
		9'd311: data = 7'd0;
		9'd312: data = 7'd11;
		9'd313: data = 7'd0;
		9'd314: data = 7'd11;
		9'd315: data = 7'd0;
		9'd316: data = 7'd11;
		9'd317: data = 7'd49;
		9'd318: data = 7'd11;
		9'd319: data = 7'd49;
		9'd320: data = 7'd0;
		9'd321: data = 7'd0;
		9'd322: data = 7'd0;
		9'd323: data = 7'd0;
		9'd324: data = 7'd2;
		9'd325: data = 7'd22;
		9'd326: data = 7'd0;
		9'd327: data = 7'd22;
		9'd328: data = 7'd21;
		9'd329: data = 7'd0;
		9'd330: data = 7'd2;
		9'd331: data = 7'd0;
		9'd332: data = 7'd0;
		9'd333: data = 7'd6;
		9'd334: data = 7'd0;
		9'd335: data = 7'd1;
		9'd336: data = 7'd1;
		9'd337: data = 7'd4;
		9'd338: data = 7'd1;
		9'd339: data = 7'd0;
		9'd340: data = 7'd2;
		9'd341: data = 7'd0;
		9'd342: data = 7'd2;
		9'd343: data = 7'd5;
		9'd344: data = 7'd2;
		9'd345: data = 7'd3;
		9'd346: data = 7'd2;
		9'd347: data = 7'd3;
		9'd348: data = 7'd21;
		9'd349: data = 7'd9;
		9'd350: data = 7'd108;
		9'd351: data = 7'd50;
		9'd352: data = 7'd3;
		9'd353: data = 7'd0;
		9'd354: data = 7'd9;
		9'd355: data = 7'd3;
		9'd356: data = 7'd0;
		9'd357: data = 7'd9;
		9'd358: data = 7'd0;
		9'd359: data = 7'd7;
		9'd360: data = 7'd0;
		9'd361: data = 7'd0;
		9'd362: data = 7'd0;
		9'd363: data = 7'd0;
		9'd364: data = 7'd109;
		9'd365: data = 7'd1;
		9'd366: data = 7'd22;
		9'd367: data = 7'd1;
		9'd368: data = 7'd0;
		9'd369: data = 7'd2;
		9'd370: data = 7'd0;
		9'd371: data = 7'd0;
		9'd372: data = 7'd0;
		9'd373: data = 7'd0;
		9'd374: data = 7'd0;
		9'd375: data = 7'd0;
		9'd376: data = 7'd0;
		9'd377: data = 7'd5;
		9'd378: data = 7'd0;
		9'd379: data = 7'd5;
		9'd380: data = 7'd0;
		9'd381: data = 7'd3;
		9'd382: data = 7'd0;
		9'd383: data = 7'd3;
		9'd384: data = 7'd5;
		9'd385: data = 7'd0;
		9'd386: data = 7'd7;
		9'd387: data = 7'd0;
		9'd388: data = 7'd0;
		9'd389: data = 7'd0;
		9'd390: data = 7'd2;
		9'd391: data = 7'd0;
		9'd392: data = 7'd0;
		9'd393: data = 7'd0;
		9'd394: data = 7'd0;
		9'd395: data = 7'd0;
		9'd396: data = 7'd0;
		9'd397: data = 7'd1;
		9'd398: data = 7'd14;
		9'd399: data = 7'd46;
		9'd400: data = 7'd0;
		9'd401: data = 7'd1;
		9'd402: data = 7'd0;
		9'd403: data = 7'd110;
		9'd404: data = 7'd0;
		9'd405: data = 7'd15;
		9'd406: data = 7'd0;
		9'd407: data = 7'd0;
		9'd408: data = 7'd0;
		9'd409: data = 7'd0;
		9'd410: data = 7'd0;
		9'd411: data = 7'd5;
		9'd412: data = 7'd0;
		9'd413: data = 7'd5;
		9'd414: data = 7'd0;
		9'd415: data = 7'd5;
		9'd416: data = 7'd0;
		9'd417: data = 7'd5;
		9'd418: data = 7'd0;
		9'd419: data = 7'd3;
		9'd420: data = 7'd0;
		9'd421: data = 7'd0;
		9'd422: data = 7'd4;
		9'd423: data = 7'd0;
		9'd424: data = 7'd0;
		9'd425: data = 7'd0;
		9'd426: data = 7'd0;
		9'd427: data = 7'd8;
		9'd428: data = 7'd0;
		9'd429: data = 7'd0;
		9'd430: data = 7'd9;
		9'd431: data = 7'd2;
		9'd432: data = 7'd22;
		9'd433: data = 7'd0;
		9'd434: data = 7'd0;
		9'd435: data = 7'd0;
		9'd436: data = 7'd0;
		9'd437: data = 7'd16;
		9'd438: data = 7'd0;
		9'd439: data = 7'd111;
		9'd440: data = 7'd0;
		9'd441: data = 7'd15;
		9'd442: data = 7'd0;
		9'd443: data = 7'd0;
		9'd444: data = 7'd0;
		9'd445: data = 7'd0;
		9'd446: data = 7'd0;
		9'd447: data = 7'd5;
		9'd448: data = 7'd0;
		9'd449: data = 7'd0;
		9'd450: data = 7'd0;
		9'd451: data = 7'd0;
		9'd452: data = 7'd8;
		9'd453: data = 7'd0;
		9'd454: data = 7'd2;
		9'd455: data = 7'd0;
		9'd456: data = 7'd0;
		9'd457: data = 7'd0;
		9'd458: data = 7'd6;
		9'd459: data = 7'd0;
		9'd460: data = 7'd0;
		9'd461: data = 7'd0;
		9'd462: data = 7'd0;
		9'd463: data = 7'd1;
		9'd464: data = 7'd7;
		9'd465: data = 7'd0;
		9'd466: data = 7'd0;
		9'd467: data = 7'd0;
		9'd468: data = 7'd0;
		9'd469: data = 7'd0;
		9'd470: data = 7'd0;
		9'd471: data = 7'd16;
		9'd472: data = 7'd0;
		9'd473: data = 7'd16;
		9'd474: data = 7'd0;
		9'd475: data = 7'd15;
		9'd476: data = 7'd0;
		9'd477: data = 7'd15;
		9'd478: data = 7'd0;
		9'd479: data = 7'd0;
		9'd480: data = 7'd0;
		9'd481: data = 7'd0;
		9'd482: data = 7'd0;
		9'd483: data = 7'd0;
		9'd484: data = 7'd4;
		9'd485: data = 7'd0;
		9'd486: data = 7'd1;
		9'd487: data = 7'd0;
		9'd488: data = 7'd6;
		9'd489: data = 7'd0;
		9'd490: data = 7'd10;
		9'd491: data = 7'd0;
		9'd492: data = 7'd0;
		9'd493: data = 7'd47;
		9'd494: data = 7'd0;
		9'd495: data = 7'd1;
		9'd496: data = 7'd0;
		9'd497: data = 7'd4;
		9'd498: data = 7'd35;
		9'd499: data = 7'd0;
		9'd500: data = 7'd0;
		9'd501: data = 7'd0;
		9'd502: data = 7'd0;
		9'd503: data = 7'd112;
		9'd504: data = 7'd0;
		9'd505: data = 7'd50;
		9'd506: data = 7'd0;
		9'd507: data = 7'd16;
		9'd508: data = 7'd0;
		9'd509: data = 7'd16;
		9'd510: data = 7'd0;
		9'd511: data = 7'd15;
		default: data = 7'd0;
	endcase
end
endmodule

module layer0_N6_rsh_1(address, data);
input wire [8:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		9'd0: data = 2'd0;
		9'd1: data = 2'd0;
		9'd2: data = 2'd1;
		9'd3: data = 2'd0;
		9'd4: data = 2'd2;
		9'd5: data = 2'd0;
		9'd6: data = 2'd2;
		9'd7: data = 2'd0;
		9'd8: data = 2'd1;
		9'd9: data = 2'd0;
		9'd10: data = 2'd2;
		9'd11: data = 2'd0;
		9'd12: data = 2'd2;
		9'd13: data = 2'd0;
		9'd14: data = 2'd0;
		9'd15: data = 2'd0;
		9'd16: data = 2'd1;
		9'd17: data = 2'd0;
		9'd18: data = 2'd2;
		9'd19: data = 2'd0;
		9'd20: data = 2'd2;
		9'd21: data = 2'd0;
		9'd22: data = 2'd2;
		9'd23: data = 2'd0;
		9'd24: data = 2'd2;
		9'd25: data = 2'd0;
		9'd26: data = 2'd0;
		9'd27: data = 2'd0;
		9'd28: data = 2'd1;
		9'd29: data = 2'd0;
		9'd30: data = 2'd2;
		9'd31: data = 2'd0;
		9'd32: data = 2'd0;
		9'd33: data = 2'd1;
		9'd34: data = 2'd0;
		9'd35: data = 2'd1;
		9'd36: data = 2'd0;
		9'd37: data = 2'd1;
		9'd38: data = 2'd0;
		9'd39: data = 2'd1;
		9'd40: data = 2'd0;
		9'd41: data = 2'd0;
		9'd42: data = 2'd0;
		9'd43: data = 2'd0;
		9'd44: data = 2'd0;
		9'd45: data = 2'd0;
		9'd46: data = 2'd0;
		9'd47: data = 2'd0;
		9'd48: data = 2'd0;
		9'd49: data = 2'd0;
		9'd50: data = 2'd0;
		9'd51: data = 2'd0;
		9'd52: data = 2'd0;
		9'd53: data = 2'd0;
		9'd54: data = 2'd0;
		9'd55: data = 2'd0;
		9'd56: data = 2'd0;
		9'd57: data = 2'd0;
		9'd58: data = 2'd2;
		9'd59: data = 2'd0;
		9'd60: data = 2'd2;
		9'd61: data = 2'd0;
		9'd62: data = 2'd0;
		9'd63: data = 2'd0;
		9'd64: data = 2'd0;
		9'd65: data = 2'd1;
		9'd66: data = 2'd0;
		9'd67: data = 2'd1;
		9'd68: data = 2'd0;
		9'd69: data = 2'd0;
		9'd70: data = 2'd0;
		9'd71: data = 2'd0;
		9'd72: data = 2'd0;
		9'd73: data = 2'd0;
		9'd74: data = 2'd0;
		9'd75: data = 2'd0;
		9'd76: data = 2'd0;
		9'd77: data = 2'd0;
		9'd78: data = 2'd0;
		9'd79: data = 2'd0;
		9'd80: data = 2'd0;
		9'd81: data = 2'd0;
		9'd82: data = 2'd0;
		9'd83: data = 2'd0;
		9'd84: data = 2'd0;
		9'd85: data = 2'd0;
		9'd86: data = 2'd0;
		9'd87: data = 2'd0;
		9'd88: data = 2'd0;
		9'd89: data = 2'd0;
		9'd90: data = 2'd0;
		9'd91: data = 2'd0;
		9'd92: data = 2'd0;
		9'd93: data = 2'd0;
		9'd94: data = 2'd0;
		9'd95: data = 2'd0;
		9'd96: data = 2'd0;
		9'd97: data = 2'd1;
		9'd98: data = 2'd0;
		9'd99: data = 2'd1;
		9'd100: data = 2'd0;
		9'd101: data = 2'd1;
		9'd102: data = 2'd0;
		9'd103: data = 2'd1;
		9'd104: data = 2'd0;
		9'd105: data = 2'd0;
		9'd106: data = 2'd0;
		9'd107: data = 2'd0;
		9'd108: data = 2'd0;
		9'd109: data = 2'd1;
		9'd110: data = 2'd0;
		9'd111: data = 2'd0;
		9'd112: data = 2'd0;
		9'd113: data = 2'd0;
		9'd114: data = 2'd0;
		9'd115: data = 2'd0;
		9'd116: data = 2'd0;
		9'd117: data = 2'd0;
		9'd118: data = 2'd0;
		9'd119: data = 2'd0;
		9'd120: data = 2'd0;
		9'd121: data = 2'd0;
		9'd122: data = 2'd0;
		9'd123: data = 2'd0;
		9'd124: data = 2'd0;
		9'd125: data = 2'd0;
		9'd126: data = 2'd0;
		9'd127: data = 2'd0;
		9'd128: data = 2'd0;
		9'd129: data = 2'd1;
		9'd130: data = 2'd0;
		9'd131: data = 2'd1;
		9'd132: data = 2'd0;
		9'd133: data = 2'd1;
		9'd134: data = 2'd0;
		9'd135: data = 2'd1;
		9'd136: data = 2'd0;
		9'd137: data = 2'd2;
		9'd138: data = 2'd0;
		9'd139: data = 2'd0;
		9'd140: data = 2'd0;
		9'd141: data = 2'd1;
		9'd142: data = 2'd0;
		9'd143: data = 2'd1;
		9'd144: data = 2'd0;
		9'd145: data = 2'd0;
		9'd146: data = 2'd0;
		9'd147: data = 2'd0;
		9'd148: data = 2'd0;
		9'd149: data = 2'd0;
		9'd150: data = 2'd0;
		9'd151: data = 2'd1;
		9'd152: data = 2'd0;
		9'd153: data = 2'd0;
		9'd154: data = 2'd0;
		9'd155: data = 2'd0;
		9'd156: data = 2'd0;
		9'd157: data = 2'd0;
		9'd158: data = 2'd0;
		9'd159: data = 2'd1;
		9'd160: data = 2'd0;
		9'd161: data = 2'd0;
		9'd162: data = 2'd0;
		9'd163: data = 2'd1;
		9'd164: data = 2'd0;
		9'd165: data = 2'd1;
		9'd166: data = 2'd0;
		9'd167: data = 2'd2;
		9'd168: data = 2'd1;
		9'd169: data = 2'd2;
		9'd170: data = 2'd1;
		9'd171: data = 2'd2;
		9'd172: data = 2'd0;
		9'd173: data = 2'd2;
		9'd174: data = 2'd0;
		9'd175: data = 2'd2;
		9'd176: data = 2'd0;
		9'd177: data = 2'd2;
		9'd178: data = 2'd0;
		9'd179: data = 2'd1;
		9'd180: data = 2'd0;
		9'd181: data = 2'd1;
		9'd182: data = 2'd0;
		9'd183: data = 2'd1;
		9'd184: data = 2'd0;
		9'd185: data = 2'd2;
		9'd186: data = 2'd0;
		9'd187: data = 2'd0;
		9'd188: data = 2'd0;
		9'd189: data = 2'd1;
		9'd190: data = 2'd0;
		9'd191: data = 2'd1;
		9'd192: data = 2'd0;
		9'd193: data = 2'd1;
		9'd194: data = 2'd0;
		9'd195: data = 2'd1;
		9'd196: data = 2'd0;
		9'd197: data = 2'd1;
		9'd198: data = 2'd0;
		9'd199: data = 2'd1;
		9'd200: data = 2'd1;
		9'd201: data = 2'd1;
		9'd202: data = 2'd2;
		9'd203: data = 2'd1;
		9'd204: data = 2'd2;
		9'd205: data = 2'd1;
		9'd206: data = 2'd2;
		9'd207: data = 2'd1;
		9'd208: data = 2'd0;
		9'd209: data = 2'd1;
		9'd210: data = 2'd0;
		9'd211: data = 2'd0;
		9'd212: data = 2'd0;
		9'd213: data = 2'd2;
		9'd214: data = 2'd0;
		9'd215: data = 2'd0;
		9'd216: data = 2'd0;
		9'd217: data = 2'd1;
		9'd218: data = 2'd0;
		9'd219: data = 2'd2;
		9'd220: data = 2'd0;
		9'd221: data = 2'd2;
		9'd222: data = 2'd0;
		9'd223: data = 2'd2;
		9'd224: data = 2'd2;
		9'd225: data = 2'd0;
		9'd226: data = 2'd2;
		9'd227: data = 2'd0;
		9'd228: data = 2'd1;
		9'd229: data = 2'd2;
		9'd230: data = 2'd0;
		9'd231: data = 2'd2;
		9'd232: data = 2'd1;
		9'd233: data = 2'd2;
		9'd234: data = 2'd1;
		9'd235: data = 2'd2;
		9'd236: data = 2'd1;
		9'd237: data = 2'd2;
		9'd238: data = 2'd1;
		9'd239: data = 2'd1;
		9'd240: data = 2'd1;
		9'd241: data = 2'd0;
		9'd242: data = 2'd0;
		9'd243: data = 2'd0;
		9'd244: data = 2'd0;
		9'd245: data = 2'd2;
		9'd246: data = 2'd0;
		9'd247: data = 2'd2;
		9'd248: data = 2'd0;
		9'd249: data = 2'd2;
		9'd250: data = 2'd0;
		9'd251: data = 2'd2;
		9'd252: data = 2'd0;
		9'd253: data = 2'd2;
		9'd254: data = 2'd0;
		9'd255: data = 2'd1;
		9'd256: data = 2'd2;
		9'd257: data = 2'd1;
		9'd258: data = 2'd1;
		9'd259: data = 2'd1;
		9'd260: data = 2'd1;
		9'd261: data = 2'd1;
		9'd262: data = 2'd1;
		9'd263: data = 2'd2;
		9'd264: data = 2'd0;
		9'd265: data = 2'd2;
		9'd266: data = 2'd1;
		9'd267: data = 2'd2;
		9'd268: data = 2'd0;
		9'd269: data = 2'd0;
		9'd270: data = 2'd1;
		9'd271: data = 2'd0;
		9'd272: data = 2'd1;
		9'd273: data = 2'd0;
		9'd274: data = 2'd1;
		9'd275: data = 2'd1;
		9'd276: data = 2'd0;
		9'd277: data = 2'd2;
		9'd278: data = 2'd0;
		9'd279: data = 2'd2;
		9'd280: data = 2'd0;
		9'd281: data = 2'd2;
		9'd282: data = 2'd0;
		9'd283: data = 2'd2;
		9'd284: data = 2'd0;
		9'd285: data = 2'd2;
		9'd286: data = 2'd0;
		9'd287: data = 2'd1;
		9'd288: data = 2'd2;
		9'd289: data = 2'd2;
		9'd290: data = 2'd2;
		9'd291: data = 2'd2;
		9'd292: data = 2'd2;
		9'd293: data = 2'd2;
		9'd294: data = 2'd0;
		9'd295: data = 2'd2;
		9'd296: data = 2'd0;
		9'd297: data = 2'd2;
		9'd298: data = 2'd1;
		9'd299: data = 2'd2;
		9'd300: data = 2'd0;
		9'd301: data = 2'd1;
		9'd302: data = 2'd0;
		9'd303: data = 2'd2;
		9'd304: data = 2'd0;
		9'd305: data = 2'd2;
		9'd306: data = 2'd1;
		9'd307: data = 2'd1;
		9'd308: data = 2'd0;
		9'd309: data = 2'd1;
		9'd310: data = 2'd0;
		9'd311: data = 2'd1;
		9'd312: data = 2'd0;
		9'd313: data = 2'd1;
		9'd314: data = 2'd0;
		9'd315: data = 2'd1;
		9'd316: data = 2'd0;
		9'd317: data = 2'd0;
		9'd318: data = 2'd0;
		9'd319: data = 2'd0;
		9'd320: data = 2'd2;
		9'd321: data = 2'd2;
		9'd322: data = 2'd1;
		9'd323: data = 2'd2;
		9'd324: data = 2'd2;
		9'd325: data = 2'd0;
		9'd326: data = 2'd0;
		9'd327: data = 2'd0;
		9'd328: data = 2'd0;
		9'd329: data = 2'd2;
		9'd330: data = 2'd2;
		9'd331: data = 2'd2;
		9'd332: data = 2'd0;
		9'd333: data = 2'd0;
		9'd334: data = 2'd1;
		9'd335: data = 2'd2;
		9'd336: data = 2'd2;
		9'd337: data = 2'd2;
		9'd338: data = 2'd2;
		9'd339: data = 2'd2;
		9'd340: data = 2'd2;
		9'd341: data = 2'd2;
		9'd342: data = 2'd2;
		9'd343: data = 2'd2;
		9'd344: data = 2'd2;
		9'd345: data = 2'd2;
		9'd346: data = 2'd2;
		9'd347: data = 2'd2;
		9'd348: data = 2'd0;
		9'd349: data = 2'd1;
		9'd350: data = 2'd0;
		9'd351: data = 2'd0;
		9'd352: data = 2'd2;
		9'd353: data = 2'd2;
		9'd354: data = 2'd1;
		9'd355: data = 2'd2;
		9'd356: data = 2'd2;
		9'd357: data = 2'd1;
		9'd358: data = 2'd2;
		9'd359: data = 2'd1;
		9'd360: data = 2'd2;
		9'd361: data = 2'd2;
		9'd362: data = 2'd2;
		9'd363: data = 2'd1;
		9'd364: data = 2'd0;
		9'd365: data = 2'd2;
		9'd366: data = 2'd0;
		9'd367: data = 2'd2;
		9'd368: data = 2'd2;
		9'd369: data = 2'd2;
		9'd370: data = 2'd2;
		9'd371: data = 2'd2;
		9'd372: data = 2'd2;
		9'd373: data = 2'd2;
		9'd374: data = 2'd2;
		9'd375: data = 2'd2;
		9'd376: data = 2'd2;
		9'd377: data = 2'd2;
		9'd378: data = 2'd2;
		9'd379: data = 2'd2;
		9'd380: data = 2'd2;
		9'd381: data = 2'd2;
		9'd382: data = 2'd2;
		9'd383: data = 2'd2;
		9'd384: data = 2'd2;
		9'd385: data = 2'd2;
		9'd386: data = 2'd1;
		9'd387: data = 2'd2;
		9'd388: data = 2'd2;
		9'd389: data = 2'd2;
		9'd390: data = 2'd2;
		9'd391: data = 2'd2;
		9'd392: data = 2'd1;
		9'd393: data = 2'd1;
		9'd394: data = 2'd2;
		9'd395: data = 2'd2;
		9'd396: data = 2'd2;
		9'd397: data = 2'd2;
		9'd398: data = 2'd1;
		9'd399: data = 2'd0;
		9'd400: data = 2'd2;
		9'd401: data = 2'd2;
		9'd402: data = 2'd2;
		9'd403: data = 2'd0;
		9'd404: data = 2'd2;
		9'd405: data = 2'd0;
		9'd406: data = 2'd2;
		9'd407: data = 2'd2;
		9'd408: data = 2'd2;
		9'd409: data = 2'd2;
		9'd410: data = 2'd2;
		9'd411: data = 2'd2;
		9'd412: data = 2'd2;
		9'd413: data = 2'd2;
		9'd414: data = 2'd2;
		9'd415: data = 2'd2;
		9'd416: data = 2'd2;
		9'd417: data = 2'd2;
		9'd418: data = 2'd2;
		9'd419: data = 2'd2;
		9'd420: data = 2'd2;
		9'd421: data = 2'd2;
		9'd422: data = 2'd2;
		9'd423: data = 2'd2;
		9'd424: data = 2'd1;
		9'd425: data = 2'd1;
		9'd426: data = 2'd2;
		9'd427: data = 2'd1;
		9'd428: data = 2'd2;
		9'd429: data = 2'd1;
		9'd430: data = 2'd1;
		9'd431: data = 2'd2;
		9'd432: data = 2'd0;
		9'd433: data = 2'd1;
		9'd434: data = 2'd2;
		9'd435: data = 2'd1;
		9'd436: data = 2'd2;
		9'd437: data = 2'd0;
		9'd438: data = 2'd2;
		9'd439: data = 2'd0;
		9'd440: data = 2'd2;
		9'd441: data = 2'd0;
		9'd442: data = 2'd2;
		9'd443: data = 2'd2;
		9'd444: data = 2'd2;
		9'd445: data = 2'd2;
		9'd446: data = 2'd2;
		9'd447: data = 2'd2;
		9'd448: data = 2'd2;
		9'd449: data = 2'd2;
		9'd450: data = 2'd2;
		9'd451: data = 2'd2;
		9'd452: data = 2'd1;
		9'd453: data = 2'd2;
		9'd454: data = 2'd2;
		9'd455: data = 2'd2;
		9'd456: data = 2'd2;
		9'd457: data = 2'd2;
		9'd458: data = 2'd0;
		9'd459: data = 2'd1;
		9'd460: data = 2'd2;
		9'd461: data = 2'd1;
		9'd462: data = 2'd2;
		9'd463: data = 2'd2;
		9'd464: data = 2'd1;
		9'd465: data = 2'd2;
		9'd466: data = 2'd2;
		9'd467: data = 2'd2;
		9'd468: data = 2'd2;
		9'd469: data = 2'd1;
		9'd470: data = 2'd2;
		9'd471: data = 2'd0;
		9'd472: data = 2'd2;
		9'd473: data = 2'd0;
		9'd474: data = 2'd2;
		9'd475: data = 2'd0;
		9'd476: data = 2'd2;
		9'd477: data = 2'd0;
		9'd478: data = 2'd2;
		9'd479: data = 2'd2;
		9'd480: data = 2'd2;
		9'd481: data = 2'd2;
		9'd482: data = 2'd2;
		9'd483: data = 2'd2;
		9'd484: data = 2'd2;
		9'd485: data = 2'd2;
		9'd486: data = 2'd2;
		9'd487: data = 2'd2;
		9'd488: data = 2'd0;
		9'd489: data = 2'd2;
		9'd490: data = 2'd1;
		9'd491: data = 2'd1;
		9'd492: data = 2'd2;
		9'd493: data = 2'd0;
		9'd494: data = 2'd2;
		9'd495: data = 2'd2;
		9'd496: data = 2'd2;
		9'd497: data = 2'd2;
		9'd498: data = 2'd0;
		9'd499: data = 2'd2;
		9'd500: data = 2'd2;
		9'd501: data = 2'd2;
		9'd502: data = 2'd2;
		9'd503: data = 2'd0;
		9'd504: data = 2'd2;
		9'd505: data = 2'd0;
		9'd506: data = 2'd2;
		9'd507: data = 2'd0;
		9'd508: data = 2'd2;
		9'd509: data = 2'd0;
		9'd510: data = 2'd2;
		9'd511: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N6(address, data);
input wire [11:0] address;
output reg [3:0] data;

wire [6:0] i; layer0_N6_idx_1 idx_1_inst(address[11:3], i);
wire [1:0] t; layer0_N6_rsh_1 rsh_1_inst(address[11:3], t);
wire [3:0] b; layer0_N6_2 layer0_N6_2_inst(address[11:3], b);
wire [2:0] u; layer0_N6_ust_1 ust_1_inst({i, address[2:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule
