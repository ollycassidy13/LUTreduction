
module layer0_N24_ust_3(address, data);
input wire [2:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		3'd0: data = 3'd0;
		3'd1: data = 3'd2;
		3'd2: data = 3'd4;
		3'd3: data = 3'd4;
		3'd4: data = 3'd4;
		3'd5: data = 3'd4;
		3'd6: data = 3'd4;
		3'd7: data = 3'd5;
		default: data = 3'd0;
	endcase
end
endmodule

module layer0_N24_rsh_3(address, data);
input wire [0:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		1'd0: data = 2'd3;
		1'd1: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N24_3(address, data);
input wire [3:0] address;
output reg [2:0] data;

wire [1:0] t; layer0_N24_rsh_3 rsh_3_inst(address[3:3], t);
wire [2:0] u; layer0_N24_ust_3 ust_3_inst(address[2:0], u);

always @(*) begin
	data = (u >> t);
end
endmodule

module layer0_N24_ust_2(address, data);
input wire [8:0] address;
output reg [3:0] data;

always @(*) begin
	case(address)
		9'd0: data = 4'd0;
		9'd1: data = 4'd2;
		9'd2: data = 4'd0;
		9'd3: data = 4'd1;
		9'd4: data = 4'd0;
		9'd5: data = 4'd1;
		9'd6: data = 4'd0;
		9'd7: data = 4'd0;
		9'd8: data = 4'd0;
		9'd9: data = 4'd0;
		9'd10: data = 4'd0;
		9'd11: data = 4'd0;
		9'd12: data = 4'd0;
		9'd13: data = 4'd0;
		9'd14: data = 4'd0;
		9'd15: data = 4'd0;
		9'd16: data = 4'd0;
		9'd17: data = 4'd0;
		9'd18: data = 4'd0;
		9'd19: data = 4'd0;
		9'd20: data = 4'd0;
		9'd21: data = 4'd0;
		9'd22: data = 4'd0;
		9'd23: data = 4'd0;
		9'd24: data = 4'd0;
		9'd25: data = 4'd0;
		9'd26: data = 4'd0;
		9'd27: data = 4'd0;
		9'd28: data = 4'd0;
		9'd29: data = 4'd0;
		9'd30: data = 4'd0;
		9'd31: data = 4'd0;
		9'd32: data = 4'd0;
		9'd33: data = 4'd6;
		9'd34: data = 4'd0;
		9'd35: data = 4'd5;
		9'd36: data = 4'd0;
		9'd37: data = 4'd4;
		9'd38: data = 4'd0;
		9'd39: data = 4'd3;
		9'd40: data = 4'd0;
		9'd41: data = 4'd3;
		9'd42: data = 4'd0;
		9'd43: data = 4'd2;
		9'd44: data = 4'd1;
		9'd45: data = 4'd2;
		9'd46: data = 4'd1;
		9'd47: data = 4'd2;
		9'd48: data = 4'd1;
		9'd49: data = 4'd2;
		9'd50: data = 4'd2;
		9'd51: data = 4'd2;
		9'd52: data = 4'd2;
		9'd53: data = 4'd2;
		9'd54: data = 4'd2;
		9'd55: data = 4'd2;
		9'd56: data = 4'd2;
		9'd57: data = 4'd2;
		9'd58: data = 4'd2;
		9'd59: data = 4'd2;
		9'd60: data = 4'd2;
		9'd61: data = 4'd2;
		9'd62: data = 4'd2;
		9'd63: data = 4'd2;
		9'd64: data = 4'd1;
		9'd65: data = 4'd8;
		9'd66: data = 4'd1;
		9'd67: data = 4'd7;
		9'd68: data = 4'd0;
		9'd69: data = 4'd7;
		9'd70: data = 4'd1;
		9'd71: data = 4'd5;
		9'd72: data = 4'd1;
		9'd73: data = 4'd4;
		9'd74: data = 4'd1;
		9'd75: data = 4'd3;
		9'd76: data = 4'd1;
		9'd77: data = 4'd2;
		9'd78: data = 4'd1;
		9'd79: data = 4'd2;
		9'd80: data = 4'd1;
		9'd81: data = 4'd2;
		9'd82: data = 4'd2;
		9'd83: data = 4'd2;
		9'd84: data = 4'd2;
		9'd85: data = 4'd2;
		9'd86: data = 4'd3;
		9'd87: data = 4'd2;
		9'd88: data = 4'd3;
		9'd89: data = 4'd3;
		9'd90: data = 4'd3;
		9'd91: data = 4'd3;
		9'd92: data = 4'd3;
		9'd93: data = 4'd3;
		9'd94: data = 4'd3;
		9'd95: data = 4'd3;
		9'd96: data = 4'd2;
		9'd97: data = 4'd8;
		9'd98: data = 4'd0;
		9'd99: data = 4'd8;
		9'd100: data = 4'd0;
		9'd101: data = 4'd7;
		9'd102: data = 4'd0;
		9'd103: data = 4'd6;
		9'd104: data = 4'd1;
		9'd105: data = 4'd6;
		9'd106: data = 4'd1;
		9'd107: data = 4'd5;
		9'd108: data = 4'd1;
		9'd109: data = 4'd3;
		9'd110: data = 4'd1;
		9'd111: data = 4'd2;
		9'd112: data = 4'd1;
		9'd113: data = 4'd2;
		9'd114: data = 4'd2;
		9'd115: data = 4'd2;
		9'd116: data = 4'd2;
		9'd117: data = 4'd3;
		9'd118: data = 4'd2;
		9'd119: data = 4'd3;
		9'd120: data = 4'd2;
		9'd121: data = 4'd3;
		9'd122: data = 4'd2;
		9'd123: data = 4'd3;
		9'd124: data = 4'd3;
		9'd125: data = 4'd3;
		9'd126: data = 4'd3;
		9'd127: data = 4'd3;
		9'd128: data = 4'd2;
		9'd129: data = 4'd10;
		9'd130: data = 4'd0;
		9'd131: data = 4'd9;
		9'd132: data = 4'd0;
		9'd133: data = 4'd9;
		9'd134: data = 4'd0;
		9'd135: data = 4'd9;
		9'd136: data = 4'd1;
		9'd137: data = 4'd8;
		9'd138: data = 4'd1;
		9'd139: data = 4'd8;
		9'd140: data = 4'd1;
		9'd141: data = 4'd7;
		9'd142: data = 4'd2;
		9'd143: data = 4'd6;
		9'd144: data = 4'd2;
		9'd145: data = 4'd4;
		9'd146: data = 4'd3;
		9'd147: data = 4'd4;
		9'd148: data = 4'd3;
		9'd149: data = 4'd4;
		9'd150: data = 4'd3;
		9'd151: data = 4'd4;
		9'd152: data = 4'd3;
		9'd153: data = 4'd4;
		9'd154: data = 4'd3;
		9'd155: data = 4'd4;
		9'd156: data = 4'd3;
		9'd157: data = 4'd4;
		9'd158: data = 4'd3;
		9'd159: data = 4'd4;
		9'd160: data = 4'd3;
		9'd161: data = 4'd11;
		9'd162: data = 4'd1;
		9'd163: data = 4'd11;
		9'd164: data = 4'd0;
		9'd165: data = 4'd11;
		9'd166: data = 4'd0;
		9'd167: data = 4'd11;
		9'd168: data = 4'd1;
		9'd169: data = 4'd10;
		9'd170: data = 4'd1;
		9'd171: data = 4'd10;
		9'd172: data = 4'd1;
		9'd173: data = 4'd10;
		9'd174: data = 4'd2;
		9'd175: data = 4'd10;
		9'd176: data = 4'd2;
		9'd177: data = 4'd8;
		9'd178: data = 4'd2;
		9'd179: data = 4'd5;
		9'd180: data = 4'd3;
		9'd181: data = 4'd6;
		9'd182: data = 4'd3;
		9'd183: data = 4'd6;
		9'd184: data = 4'd3;
		9'd185: data = 4'd6;
		9'd186: data = 4'd3;
		9'd187: data = 4'd5;
		9'd188: data = 4'd3;
		9'd189: data = 4'd5;
		9'd190: data = 4'd3;
		9'd191: data = 4'd5;
		9'd192: data = 4'd4;
		9'd193: data = 4'd11;
		9'd194: data = 4'd1;
		9'd195: data = 4'd11;
		9'd196: data = 4'd0;
		9'd197: data = 4'd11;
		9'd198: data = 4'd0;
		9'd199: data = 4'd11;
		9'd200: data = 4'd0;
		9'd201: data = 4'd11;
		9'd202: data = 4'd1;
		9'd203: data = 4'd11;
		9'd204: data = 4'd1;
		9'd205: data = 4'd11;
		9'd206: data = 4'd2;
		9'd207: data = 4'd11;
		9'd208: data = 4'd2;
		9'd209: data = 4'd11;
		9'd210: data = 4'd2;
		9'd211: data = 4'd10;
		9'd212: data = 4'd3;
		9'd213: data = 4'd7;
		9'd214: data = 4'd3;
		9'd215: data = 4'd7;
		9'd216: data = 4'd3;
		9'd217: data = 4'd7;
		9'd218: data = 4'd3;
		9'd219: data = 4'd7;
		9'd220: data = 4'd4;
		9'd221: data = 4'd7;
		9'd222: data = 4'd4;
		9'd223: data = 4'd6;
		9'd224: data = 4'd5;
		9'd225: data = 4'd11;
		9'd226: data = 4'd2;
		9'd227: data = 4'd11;
		9'd228: data = 4'd0;
		9'd229: data = 4'd11;
		9'd230: data = 4'd0;
		9'd231: data = 4'd11;
		9'd232: data = 4'd0;
		9'd233: data = 4'd11;
		9'd234: data = 4'd0;
		9'd235: data = 4'd11;
		9'd236: data = 4'd1;
		9'd237: data = 4'd11;
		9'd238: data = 4'd2;
		9'd239: data = 4'd11;
		9'd240: data = 4'd2;
		9'd241: data = 4'd11;
		9'd242: data = 4'd2;
		9'd243: data = 4'd11;
		9'd244: data = 4'd3;
		9'd245: data = 4'd10;
		9'd246: data = 4'd3;
		9'd247: data = 4'd8;
		9'd248: data = 4'd3;
		9'd249: data = 4'd8;
		9'd250: data = 4'd4;
		9'd251: data = 4'd8;
		9'd252: data = 4'd4;
		9'd253: data = 4'd8;
		9'd254: data = 4'd5;
		9'd255: data = 4'd8;
		9'd256: data = 4'd6;
		9'd257: data = 4'd10;
		9'd258: data = 4'd4;
		9'd259: data = 4'd10;
		9'd260: data = 4'd1;
		9'd261: data = 4'd10;
		9'd262: data = 4'd0;
		9'd263: data = 4'd10;
		9'd264: data = 4'd0;
		9'd265: data = 4'd10;
		9'd266: data = 4'd0;
		9'd267: data = 4'd10;
		9'd268: data = 4'd0;
		9'd269: data = 4'd10;
		9'd270: data = 4'd1;
		9'd271: data = 4'd10;
		9'd272: data = 4'd2;
		9'd273: data = 4'd10;
		9'd274: data = 4'd2;
		9'd275: data = 4'd10;
		9'd276: data = 4'd2;
		9'd277: data = 4'd10;
		9'd278: data = 4'd3;
		9'd279: data = 4'd8;
		9'd280: data = 4'd3;
		9'd281: data = 4'd8;
		9'd282: data = 4'd4;
		9'd283: data = 4'd8;
		9'd284: data = 4'd4;
		9'd285: data = 4'd8;
		9'd286: data = 4'd4;
		9'd287: data = 4'd8;
		default: data = 4'd0;
	endcase
end
endmodule

module layer0_N24_idx_2(address, data);
input wire [3:0] address;
output reg [3:0] data;

always @(*) begin
	case(address)
		4'd0: data = 4'd0;
		4'd1: data = 4'd0;
		4'd2: data = 4'd0;
		4'd3: data = 4'd0;
		4'd4: data = 4'd0;
		4'd5: data = 4'd0;
		4'd6: data = 4'd0;
		4'd7: data = 4'd0;
		4'd8: data = 4'd1;
		4'd9: data = 4'd2;
		4'd10: data = 4'd3;
		4'd11: data = 4'd4;
		4'd12: data = 4'd5;
		4'd13: data = 4'd6;
		4'd14: data = 4'd7;
		4'd15: data = 4'd8;
		default: data = 4'd0;
	endcase
end
endmodule

module layer0_N24_rsh_2(address, data);
input wire [3:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		4'd0: data = 2'd2;
		4'd1: data = 2'd2;
		4'd2: data = 2'd2;
		4'd3: data = 2'd2;
		4'd4: data = 2'd2;
		4'd5: data = 2'd2;
		4'd6: data = 2'd2;
		4'd7: data = 2'd0;
		4'd8: data = 2'd0;
		4'd9: data = 2'd0;
		4'd10: data = 2'd0;
		4'd11: data = 2'd0;
		4'd12: data = 2'd0;
		4'd13: data = 2'd0;
		4'd14: data = 2'd0;
		4'd15: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N24_2(address, data);
input wire [8:0] address;
output reg [3:0] data;

wire [3:0] i; layer0_N24_idx_2 idx_2_inst(address[8:5], i);
wire [1:0] t; layer0_N24_rsh_2 rsh_2_inst(address[8:5], t);
wire [2:0] b; layer0_N24_3 layer0_N24_3_inst(address[8:5], b);
wire [3:0] u; layer0_N24_ust_2 ust_2_inst({i, address[4:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule

module layer0_N24_ust_1(address, data);
input wire [10:0] address;
output reg [3:0] data;

always @(*) begin
	case(address)
		11'd0: data = 4'd0;
		11'd1: data = 4'd0;
		11'd2: data = 4'd0;
		11'd3: data = 4'd0;
		11'd4: data = 4'd0;
		11'd5: data = 4'd1;
		11'd6: data = 4'd3;
		11'd7: data = 4'd4;
		11'd8: data = 4'd4;
		11'd9: data = 4'd3;
		11'd10: data = 4'd2;
		11'd11: data = 4'd1;
		11'd12: data = 4'd0;
		11'd13: data = 4'd0;
		11'd14: data = 4'd0;
		11'd15: data = 4'd0;
		11'd16: data = 4'd0;
		11'd17: data = 4'd4;
		11'd18: data = 4'd6;
		11'd19: data = 4'd6;
		11'd20: data = 4'd6;
		11'd21: data = 4'd6;
		11'd22: data = 4'd6;
		11'd23: data = 4'd6;
		11'd24: data = 4'd3;
		11'd25: data = 4'd2;
		11'd26: data = 4'd1;
		11'd27: data = 4'd0;
		11'd28: data = 4'd0;
		11'd29: data = 4'd0;
		11'd30: data = 4'd0;
		11'd31: data = 4'd0;
		11'd32: data = 4'd0;
		11'd33: data = 4'd0;
		11'd34: data = 4'd0;
		11'd35: data = 4'd0;
		11'd36: data = 4'd1;
		11'd37: data = 4'd3;
		11'd38: data = 4'd4;
		11'd39: data = 4'd6;
		11'd40: data = 4'd2;
		11'd41: data = 4'd1;
		11'd42: data = 4'd0;
		11'd43: data = 4'd0;
		11'd44: data = 4'd0;
		11'd45: data = 4'd0;
		11'd46: data = 4'd0;
		11'd47: data = 4'd0;
		11'd48: data = 4'd0;
		11'd49: data = 4'd3;
		11'd50: data = 4'd4;
		11'd51: data = 4'd4;
		11'd52: data = 4'd4;
		11'd53: data = 4'd4;
		11'd54: data = 4'd4;
		11'd55: data = 4'd4;
		11'd56: data = 4'd0;
		11'd57: data = 4'd0;
		11'd58: data = 4'd0;
		11'd59: data = 4'd1;
		11'd60: data = 4'd2;
		11'd61: data = 4'd4;
		11'd62: data = 4'd7;
		11'd63: data = 4'd9;
		11'd64: data = 4'd0;
		11'd65: data = 4'd0;
		11'd66: data = 4'd1;
		11'd67: data = 4'd2;
		11'd68: data = 4'd3;
		11'd69: data = 4'd4;
		11'd70: data = 4'd5;
		11'd71: data = 4'd6;
		11'd72: data = 4'd0;
		11'd73: data = 4'd0;
		11'd74: data = 4'd0;
		11'd75: data = 4'd0;
		11'd76: data = 4'd0;
		11'd77: data = 4'd0;
		11'd78: data = 4'd1;
		11'd79: data = 4'd4;
		11'd80: data = 4'd0;
		11'd81: data = 4'd0;
		11'd82: data = 4'd0;
		11'd83: data = 4'd0;
		11'd84: data = 4'd0;
		11'd85: data = 4'd1;
		11'd86: data = 4'd4;
		11'd87: data = 4'd7;
		11'd88: data = 4'd0;
		11'd89: data = 4'd1;
		11'd90: data = 4'd3;
		11'd91: data = 4'd4;
		11'd92: data = 4'd5;
		11'd93: data = 4'd7;
		11'd94: data = 4'd8;
		11'd95: data = 4'd10;
		11'd96: data = 4'd0;
		11'd97: data = 4'd0;
		11'd98: data = 4'd0;
		11'd99: data = 4'd1;
		11'd100: data = 4'd3;
		11'd101: data = 4'd6;
		11'd102: data = 4'd8;
		11'd103: data = 4'd10;
		11'd104: data = 4'd0;
		11'd105: data = 4'd0;
		11'd106: data = 4'd0;
		11'd107: data = 4'd0;
		11'd108: data = 4'd2;
		11'd109: data = 4'd3;
		11'd110: data = 4'd4;
		11'd111: data = 4'd5;
		11'd112: data = 4'd0;
		11'd113: data = 4'd3;
		11'd114: data = 4'd4;
		11'd115: data = 4'd4;
		11'd116: data = 4'd6;
		11'd117: data = 4'd6;
		11'd118: data = 4'd7;
		11'd119: data = 4'd7;
		11'd120: data = 4'd0;
		11'd121: data = 4'd3;
		11'd122: data = 4'd5;
		11'd123: data = 4'd6;
		11'd124: data = 4'd7;
		11'd125: data = 4'd7;
		11'd126: data = 4'd7;
		11'd127: data = 4'd7;
		11'd128: data = 4'd0;
		11'd129: data = 4'd0;
		11'd130: data = 4'd0;
		11'd131: data = 4'd0;
		11'd132: data = 4'd1;
		11'd133: data = 4'd3;
		11'd134: data = 4'd5;
		11'd135: data = 4'd8;
		11'd136: data = 4'd0;
		11'd137: data = 4'd0;
		11'd138: data = 4'd0;
		11'd139: data = 4'd0;
		11'd140: data = 4'd0;
		11'd141: data = 4'd2;
		11'd142: data = 4'd3;
		11'd143: data = 4'd4;
		11'd144: data = 4'd0;
		11'd145: data = 4'd0;
		11'd146: data = 4'd0;
		11'd147: data = 4'd2;
		11'd148: data = 4'd5;
		11'd149: data = 4'd7;
		11'd150: data = 4'd9;
		11'd151: data = 4'd11;
		11'd152: data = 4'd0;
		11'd153: data = 4'd1;
		11'd154: data = 4'd2;
		11'd155: data = 4'd5;
		11'd156: data = 4'd7;
		11'd157: data = 4'd8;
		11'd158: data = 4'd10;
		11'd159: data = 4'd11;
		11'd160: data = 4'd0;
		11'd161: data = 4'd1;
		11'd162: data = 4'd2;
		11'd163: data = 4'd4;
		11'd164: data = 4'd5;
		11'd165: data = 4'd6;
		11'd166: data = 4'd8;
		11'd167: data = 4'd9;
		11'd168: data = 4'd2;
		11'd169: data = 4'd1;
		11'd170: data = 4'd1;
		11'd171: data = 4'd1;
		11'd172: data = 4'd1;
		11'd173: data = 4'd0;
		11'd174: data = 4'd0;
		11'd175: data = 4'd0;
		11'd176: data = 4'd5;
		11'd177: data = 4'd4;
		11'd178: data = 4'd3;
		11'd179: data = 4'd2;
		11'd180: data = 4'd1;
		11'd181: data = 4'd0;
		11'd182: data = 4'd0;
		11'd183: data = 4'd0;
		11'd184: data = 4'd0;
		11'd185: data = 4'd1;
		11'd186: data = 4'd2;
		11'd187: data = 4'd3;
		11'd188: data = 4'd4;
		11'd189: data = 4'd4;
		11'd190: data = 4'd5;
		11'd191: data = 4'd5;
		11'd192: data = 4'd4;
		11'd193: data = 4'd3;
		11'd194: data = 4'd2;
		11'd195: data = 4'd1;
		11'd196: data = 4'd0;
		11'd197: data = 4'd0;
		11'd198: data = 4'd1;
		11'd199: data = 4'd2;
		11'd200: data = 4'd0;
		11'd201: data = 4'd1;
		11'd202: data = 4'd5;
		11'd203: data = 4'd9;
		11'd204: data = 4'd11;
		11'd205: data = 4'd11;
		11'd206: data = 4'd11;
		11'd207: data = 4'd11;
		11'd208: data = 4'd0;
		11'd209: data = 4'd0;
		11'd210: data = 4'd0;
		11'd211: data = 4'd0;
		11'd212: data = 4'd0;
		11'd213: data = 4'd0;
		11'd214: data = 4'd1;
		11'd215: data = 4'd3;
		11'd216: data = 4'd0;
		11'd217: data = 4'd0;
		11'd218: data = 4'd0;
		11'd219: data = 4'd0;
		11'd220: data = 4'd2;
		11'd221: data = 4'd4;
		11'd222: data = 4'd7;
		11'd223: data = 4'd10;
		11'd224: data = 4'd0;
		11'd225: data = 4'd0;
		11'd226: data = 4'd0;
		11'd227: data = 4'd0;
		11'd228: data = 4'd1;
		11'd229: data = 4'd2;
		11'd230: data = 4'd4;
		11'd231: data = 4'd5;
		11'd232: data = 4'd0;
		11'd233: data = 4'd0;
		11'd234: data = 4'd1;
		11'd235: data = 4'd2;
		11'd236: data = 4'd4;
		11'd237: data = 4'd5;
		11'd238: data = 4'd7;
		11'd239: data = 4'd9;
		11'd240: data = 4'd0;
		11'd241: data = 4'd1;
		11'd242: data = 4'd2;
		11'd243: data = 4'd4;
		11'd244: data = 4'd6;
		11'd245: data = 4'd7;
		11'd246: data = 4'd8;
		11'd247: data = 4'd10;
		11'd248: data = 4'd0;
		11'd249: data = 4'd1;
		11'd250: data = 4'd3;
		11'd251: data = 4'd4;
		11'd252: data = 4'd6;
		11'd253: data = 4'd7;
		11'd254: data = 4'd8;
		11'd255: data = 4'd9;
		11'd256: data = 4'd0;
		11'd257: data = 4'd1;
		11'd258: data = 4'd1;
		11'd259: data = 4'd2;
		11'd260: data = 4'd3;
		11'd261: data = 4'd4;
		11'd262: data = 4'd5;
		11'd263: data = 4'd6;
		11'd264: data = 4'd0;
		11'd265: data = 4'd2;
		11'd266: data = 4'd3;
		11'd267: data = 4'd4;
		11'd268: data = 4'd5;
		11'd269: data = 4'd6;
		11'd270: data = 4'd7;
		11'd271: data = 4'd8;
		11'd272: data = 4'd0;
		11'd273: data = 4'd2;
		11'd274: data = 4'd3;
		11'd275: data = 4'd4;
		11'd276: data = 4'd5;
		11'd277: data = 4'd6;
		11'd278: data = 4'd8;
		11'd279: data = 4'd9;
		11'd280: data = 4'd0;
		11'd281: data = 4'd1;
		11'd282: data = 4'd2;
		11'd283: data = 4'd2;
		11'd284: data = 4'd3;
		11'd285: data = 4'd4;
		11'd286: data = 4'd5;
		11'd287: data = 4'd5;
		11'd288: data = 4'd0;
		11'd289: data = 4'd1;
		11'd290: data = 4'd2;
		11'd291: data = 4'd3;
		11'd292: data = 4'd6;
		11'd293: data = 4'd7;
		11'd294: data = 4'd8;
		11'd295: data = 4'd9;
		11'd296: data = 4'd0;
		11'd297: data = 4'd1;
		11'd298: data = 4'd1;
		11'd299: data = 4'd2;
		11'd300: data = 4'd3;
		11'd301: data = 4'd3;
		11'd302: data = 4'd4;
		11'd303: data = 4'd5;
		11'd304: data = 4'd0;
		11'd305: data = 4'd2;
		11'd306: data = 4'd3;
		11'd307: data = 4'd4;
		11'd308: data = 4'd5;
		11'd309: data = 4'd5;
		11'd310: data = 4'd5;
		11'd311: data = 4'd5;
		11'd312: data = 4'd0;
		11'd313: data = 4'd1;
		11'd314: data = 4'd2;
		11'd315: data = 4'd2;
		11'd316: data = 4'd3;
		11'd317: data = 4'd4;
		11'd318: data = 4'd4;
		11'd319: data = 4'd5;
		11'd320: data = 4'd0;
		11'd321: data = 4'd1;
		11'd322: data = 4'd2;
		11'd323: data = 4'd3;
		11'd324: data = 4'd3;
		11'd325: data = 4'd4;
		11'd326: data = 4'd5;
		11'd327: data = 4'd5;
		11'd328: data = 4'd4;
		11'd329: data = 4'd2;
		11'd330: data = 4'd1;
		11'd331: data = 4'd0;
		11'd332: data = 4'd0;
		11'd333: data = 4'd1;
		11'd334: data = 4'd2;
		11'd335: data = 4'd3;
		11'd336: data = 4'd1;
		11'd337: data = 4'd0;
		11'd338: data = 4'd2;
		11'd339: data = 4'd5;
		11'd340: data = 4'd9;
		11'd341: data = 4'd11;
		11'd342: data = 4'd11;
		11'd343: data = 4'd11;
		11'd344: data = 4'd4;
		11'd345: data = 4'd3;
		11'd346: data = 4'd2;
		11'd347: data = 4'd1;
		11'd348: data = 4'd0;
		11'd349: data = 4'd1;
		11'd350: data = 4'd2;
		11'd351: data = 4'd3;
		11'd352: data = 4'd0;
		11'd353: data = 4'd0;
		11'd354: data = 4'd0;
		11'd355: data = 4'd0;
		11'd356: data = 4'd0;
		11'd357: data = 4'd1;
		11'd358: data = 4'd2;
		11'd359: data = 4'd5;
		11'd360: data = 4'd0;
		11'd361: data = 4'd0;
		11'd362: data = 4'd0;
		11'd363: data = 4'd0;
		11'd364: data = 4'd1;
		11'd365: data = 4'd2;
		11'd366: data = 4'd3;
		11'd367: data = 4'd6;
		11'd368: data = 4'd0;
		11'd369: data = 4'd0;
		11'd370: data = 4'd0;
		11'd371: data = 4'd0;
		11'd372: data = 4'd2;
		11'd373: data = 4'd3;
		11'd374: data = 4'd5;
		11'd375: data = 4'd8;
		11'd376: data = 4'd0;
		11'd377: data = 4'd0;
		11'd378: data = 4'd2;
		11'd379: data = 4'd3;
		11'd380: data = 4'd6;
		11'd381: data = 4'd7;
		11'd382: data = 4'd9;
		11'd383: data = 4'd10;
		11'd384: data = 4'd0;
		11'd385: data = 4'd0;
		11'd386: data = 4'd1;
		11'd387: data = 4'd3;
		11'd388: data = 4'd4;
		11'd389: data = 4'd6;
		11'd390: data = 4'd8;
		11'd391: data = 4'd9;
		11'd392: data = 4'd0;
		11'd393: data = 4'd0;
		11'd394: data = 4'd0;
		11'd395: data = 4'd2;
		11'd396: data = 4'd3;
		11'd397: data = 4'd5;
		11'd398: data = 4'd6;
		11'd399: data = 4'd8;
		11'd400: data = 4'd0;
		11'd401: data = 4'd0;
		11'd402: data = 4'd0;
		11'd403: data = 4'd1;
		11'd404: data = 4'd3;
		11'd405: data = 4'd4;
		11'd406: data = 4'd5;
		11'd407: data = 4'd7;
		11'd408: data = 4'd0;
		11'd409: data = 4'd0;
		11'd410: data = 4'd0;
		11'd411: data = 4'd1;
		11'd412: data = 4'd2;
		11'd413: data = 4'd3;
		11'd414: data = 4'd5;
		11'd415: data = 4'd6;
		11'd416: data = 4'd0;
		11'd417: data = 4'd1;
		11'd418: data = 4'd2;
		11'd419: data = 4'd4;
		11'd420: data = 4'd5;
		11'd421: data = 4'd7;
		11'd422: data = 4'd8;
		11'd423: data = 4'd9;
		11'd424: data = 4'd0;
		11'd425: data = 4'd0;
		11'd426: data = 4'd2;
		11'd427: data = 4'd3;
		11'd428: data = 4'd4;
		11'd429: data = 4'd6;
		11'd430: data = 4'd8;
		11'd431: data = 4'd9;
		11'd432: data = 4'd0;
		11'd433: data = 4'd0;
		11'd434: data = 4'd1;
		11'd435: data = 4'd2;
		11'd436: data = 4'd3;
		11'd437: data = 4'd4;
		11'd438: data = 4'd6;
		11'd439: data = 4'd8;
		11'd440: data = 4'd0;
		11'd441: data = 4'd0;
		11'd442: data = 4'd1;
		11'd443: data = 4'd2;
		11'd444: data = 4'd3;
		11'd445: data = 4'd4;
		11'd446: data = 4'd5;
		11'd447: data = 4'd7;
		11'd448: data = 4'd0;
		11'd449: data = 4'd0;
		11'd450: data = 4'd1;
		11'd451: data = 4'd1;
		11'd452: data = 4'd2;
		11'd453: data = 4'd4;
		11'd454: data = 4'd5;
		11'd455: data = 4'd6;
		11'd456: data = 4'd5;
		11'd457: data = 4'd4;
		11'd458: data = 4'd3;
		11'd459: data = 4'd2;
		11'd460: data = 4'd0;
		11'd461: data = 4'd0;
		11'd462: data = 4'd0;
		11'd463: data = 4'd0;
		11'd464: data = 4'd0;
		11'd465: data = 4'd0;
		11'd466: data = 4'd0;
		11'd467: data = 4'd1;
		11'd468: data = 4'd2;
		11'd469: data = 4'd4;
		11'd470: data = 4'd5;
		11'd471: data = 4'd6;
		11'd472: data = 4'd0;
		11'd473: data = 4'd0;
		11'd474: data = 4'd0;
		11'd475: data = 4'd0;
		11'd476: data = 4'd1;
		11'd477: data = 4'd2;
		11'd478: data = 4'd2;
		11'd479: data = 4'd4;
		11'd480: data = 4'd1;
		11'd481: data = 4'd1;
		11'd482: data = 4'd0;
		11'd483: data = 4'd0;
		11'd484: data = 4'd0;
		11'd485: data = 4'd1;
		11'd486: data = 4'd1;
		11'd487: data = 4'd2;
		11'd488: data = 4'd0;
		11'd489: data = 4'd1;
		11'd490: data = 4'd3;
		11'd491: data = 4'd4;
		11'd492: data = 4'd6;
		11'd493: data = 4'd7;
		11'd494: data = 4'd8;
		11'd495: data = 4'd10;
		11'd496: data = 4'd2;
		11'd497: data = 4'd1;
		11'd498: data = 4'd1;
		11'd499: data = 4'd1;
		11'd500: data = 4'd0;
		11'd501: data = 4'd0;
		11'd502: data = 4'd1;
		11'd503: data = 4'd2;
		11'd504: data = 4'd3;
		11'd505: data = 4'd2;
		11'd506: data = 4'd2;
		11'd507: data = 4'd1;
		11'd508: data = 4'd1;
		11'd509: data = 4'd0;
		11'd510: data = 4'd1;
		11'd511: data = 4'd1;
		11'd512: data = 4'd0;
		11'd513: data = 4'd1;
		11'd514: data = 4'd2;
		11'd515: data = 4'd4;
		11'd516: data = 4'd5;
		11'd517: data = 4'd7;
		11'd518: data = 4'd8;
		11'd519: data = 4'd10;
		11'd520: data = 4'd2;
		11'd521: data = 4'd1;
		11'd522: data = 4'd1;
		11'd523: data = 4'd1;
		11'd524: data = 4'd0;
		11'd525: data = 4'd0;
		11'd526: data = 4'd0;
		11'd527: data = 4'd0;
		11'd528: data = 4'd0;
		11'd529: data = 4'd1;
		11'd530: data = 4'd2;
		11'd531: data = 4'd3;
		11'd532: data = 4'd5;
		11'd533: data = 4'd6;
		11'd534: data = 4'd8;
		11'd535: data = 4'd9;
		11'd536: data = 4'd0;
		11'd537: data = 4'd0;
		11'd538: data = 4'd1;
		11'd539: data = 4'd2;
		11'd540: data = 4'd3;
		11'd541: data = 4'd6;
		11'd542: data = 4'd7;
		11'd543: data = 4'd9;
		11'd544: data = 4'd3;
		11'd545: data = 4'd2;
		11'd546: data = 4'd1;
		11'd547: data = 4'd1;
		11'd548: data = 4'd1;
		11'd549: data = 4'd1;
		11'd550: data = 4'd0;
		11'd551: data = 4'd0;
		11'd552: data = 4'd0;
		11'd553: data = 4'd0;
		11'd554: data = 4'd1;
		11'd555: data = 4'd2;
		11'd556: data = 4'd3;
		11'd557: data = 4'd5;
		11'd558: data = 4'd7;
		11'd559: data = 4'd8;
		11'd560: data = 4'd0;
		11'd561: data = 4'd0;
		11'd562: data = 4'd1;
		11'd563: data = 4'd2;
		11'd564: data = 4'd3;
		11'd565: data = 4'd4;
		11'd566: data = 4'd5;
		11'd567: data = 4'd8;
		11'd568: data = 4'd0;
		11'd569: data = 4'd1;
		11'd570: data = 4'd1;
		11'd571: data = 4'd2;
		11'd572: data = 4'd3;
		11'd573: data = 4'd4;
		11'd574: data = 4'd5;
		11'd575: data = 4'd5;
		11'd576: data = 4'd0;
		11'd577: data = 4'd0;
		11'd578: data = 4'd0;
		11'd579: data = 4'd1;
		11'd580: data = 4'd1;
		11'd581: data = 4'd2;
		11'd582: data = 4'd5;
		11'd583: data = 4'd6;
		11'd584: data = 4'd0;
		11'd585: data = 4'd0;
		11'd586: data = 4'd0;
		11'd587: data = 4'd0;
		11'd588: data = 4'd0;
		11'd589: data = 4'd1;
		11'd590: data = 4'd3;
		11'd591: data = 4'd5;
		11'd592: data = 4'd0;
		11'd593: data = 4'd1;
		11'd594: data = 4'd2;
		11'd595: data = 4'd3;
		11'd596: data = 4'd4;
		11'd597: data = 4'd4;
		11'd598: data = 4'd5;
		11'd599: data = 4'd6;
		11'd600: data = 4'd0;
		11'd601: data = 4'd1;
		11'd602: data = 4'd1;
		11'd603: data = 4'd1;
		11'd604: data = 4'd1;
		11'd605: data = 4'd1;
		11'd606: data = 4'd2;
		11'd607: data = 4'd4;
		11'd608: data = 4'd0;
		11'd609: data = 4'd2;
		11'd610: data = 4'd3;
		11'd611: data = 4'd4;
		11'd612: data = 4'd5;
		11'd613: data = 4'd6;
		11'd614: data = 4'd6;
		11'd615: data = 4'd7;
		11'd616: data = 4'd1;
		11'd617: data = 4'd1;
		11'd618: data = 4'd1;
		11'd619: data = 4'd0;
		11'd620: data = 4'd0;
		11'd621: data = 4'd0;
		11'd622: data = 4'd0;
		11'd623: data = 4'd1;
		11'd624: data = 4'd0;
		11'd625: data = 4'd2;
		11'd626: data = 4'd4;
		11'd627: data = 4'd5;
		11'd628: data = 4'd6;
		11'd629: data = 4'd6;
		11'd630: data = 4'd7;
		11'd631: data = 4'd8;
		11'd632: data = 4'd2;
		11'd633: data = 4'd1;
		11'd634: data = 4'd1;
		11'd635: data = 4'd1;
		11'd636: data = 4'd0;
		11'd637: data = 4'd0;
		11'd638: data = 4'd0;
		11'd639: data = 4'd1;
		11'd640: data = 4'd0;
		11'd641: data = 4'd2;
		11'd642: data = 4'd4;
		11'd643: data = 4'd5;
		11'd644: data = 4'd6;
		11'd645: data = 4'd7;
		11'd646: data = 4'd8;
		11'd647: data = 4'd9;
		11'd648: data = 4'd0;
		11'd649: data = 4'd1;
		11'd650: data = 4'd4;
		11'd651: data = 4'd6;
		11'd652: data = 4'd7;
		11'd653: data = 4'd8;
		11'd654: data = 4'd9;
		11'd655: data = 4'd10;
		11'd656: data = 4'd3;
		11'd657: data = 4'd2;
		11'd658: data = 4'd2;
		11'd659: data = 4'd1;
		11'd660: data = 4'd1;
		11'd661: data = 4'd1;
		11'd662: data = 4'd0;
		11'd663: data = 4'd0;
		11'd664: data = 4'd0;
		11'd665: data = 4'd1;
		11'd666: data = 4'd2;
		11'd667: data = 4'd5;
		11'd668: data = 4'd7;
		11'd669: data = 4'd8;
		11'd670: data = 4'd9;
		11'd671: data = 4'd9;
		11'd672: data = 4'd3;
		11'd673: data = 4'd2;
		11'd674: data = 4'd2;
		11'd675: data = 4'd2;
		11'd676: data = 4'd1;
		11'd677: data = 4'd1;
		11'd678: data = 4'd1;
		11'd679: data = 4'd0;
		11'd680: data = 4'd2;
		11'd681: data = 4'd2;
		11'd682: data = 4'd1;
		11'd683: data = 4'd1;
		11'd684: data = 4'd1;
		11'd685: data = 4'd1;
		11'd686: data = 4'd0;
		11'd687: data = 4'd0;
		11'd688: data = 4'd0;
		11'd689: data = 4'd1;
		11'd690: data = 4'd2;
		11'd691: data = 4'd3;
		11'd692: data = 4'd3;
		11'd693: data = 4'd6;
		11'd694: data = 4'd8;
		11'd695: data = 4'd9;
		11'd696: data = 4'd3;
		11'd697: data = 4'd2;
		11'd698: data = 4'd1;
		11'd699: data = 4'd1;
		11'd700: data = 4'd1;
		11'd701: data = 4'd1;
		11'd702: data = 4'd1;
		11'd703: data = 4'd0;
		11'd704: data = 4'd0;
		11'd705: data = 4'd1;
		11'd706: data = 4'd2;
		11'd707: data = 4'd3;
		11'd708: data = 4'd3;
		11'd709: data = 4'd4;
		11'd710: data = 4'd6;
		11'd711: data = 4'd8;
		11'd712: data = 4'd0;
		11'd713: data = 4'd1;
		11'd714: data = 4'd2;
		11'd715: data = 4'd3;
		11'd716: data = 4'd3;
		11'd717: data = 4'd4;
		11'd718: data = 4'd5;
		11'd719: data = 4'd6;
		11'd720: data = 4'd3;
		11'd721: data = 4'd3;
		11'd722: data = 4'd2;
		11'd723: data = 4'd1;
		11'd724: data = 4'd0;
		11'd725: data = 4'd0;
		11'd726: data = 4'd0;
		11'd727: data = 4'd0;
		11'd728: data = 4'd0;
		11'd729: data = 4'd1;
		11'd730: data = 4'd1;
		11'd731: data = 4'd2;
		11'd732: data = 4'd2;
		11'd733: data = 4'd4;
		11'd734: data = 4'd4;
		11'd735: data = 4'd5;
		11'd736: data = 4'd0;
		11'd737: data = 4'd2;
		11'd738: data = 4'd2;
		11'd739: data = 4'd2;
		11'd740: data = 4'd2;
		11'd741: data = 4'd4;
		11'd742: data = 4'd6;
		11'd743: data = 4'd7;
		11'd744: data = 4'd0;
		11'd745: data = 4'd0;
		11'd746: data = 4'd1;
		11'd747: data = 4'd2;
		11'd748: data = 4'd2;
		11'd749: data = 4'd3;
		11'd750: data = 4'd3;
		11'd751: data = 4'd3;
		11'd752: data = 4'd0;
		11'd753: data = 4'd1;
		11'd754: data = 4'd1;
		11'd755: data = 4'd1;
		11'd756: data = 4'd1;
		11'd757: data = 4'd2;
		11'd758: data = 4'd4;
		11'd759: data = 4'd6;
		11'd760: data = 4'd0;
		11'd761: data = 4'd1;
		11'd762: data = 4'd1;
		11'd763: data = 4'd2;
		11'd764: data = 4'd3;
		11'd765: data = 4'd4;
		11'd766: data = 4'd4;
		11'd767: data = 4'd4;
		11'd768: data = 4'd0;
		11'd769: data = 4'd0;
		11'd770: data = 4'd1;
		11'd771: data = 4'd1;
		11'd772: data = 4'd1;
		11'd773: data = 4'd1;
		11'd774: data = 4'd3;
		11'd775: data = 4'd5;
		11'd776: data = 4'd0;
		11'd777: data = 4'd1;
		11'd778: data = 4'd2;
		11'd779: data = 4'd3;
		11'd780: data = 4'd4;
		11'd781: data = 4'd5;
		11'd782: data = 4'd5;
		11'd783: data = 4'd5;
		11'd784: data = 4'd0;
		11'd785: data = 4'd0;
		11'd786: data = 4'd0;
		11'd787: data = 4'd0;
		11'd788: data = 4'd0;
		11'd789: data = 4'd0;
		11'd790: data = 4'd0;
		11'd791: data = 4'd3;
		11'd792: data = 4'd1;
		11'd793: data = 4'd0;
		11'd794: data = 4'd1;
		11'd795: data = 4'd1;
		11'd796: data = 4'd0;
		11'd797: data = 4'd0;
		11'd798: data = 4'd0;
		11'd799: data = 4'd1;
		11'd800: data = 4'd0;
		11'd801: data = 4'd2;
		11'd802: data = 4'd3;
		11'd803: data = 4'd4;
		11'd804: data = 4'd4;
		11'd805: data = 4'd5;
		11'd806: data = 4'd6;
		11'd807: data = 4'd6;
		11'd808: data = 4'd0;
		11'd809: data = 4'd3;
		11'd810: data = 4'd4;
		11'd811: data = 4'd5;
		11'd812: data = 4'd6;
		11'd813: data = 4'd7;
		11'd814: data = 4'd8;
		11'd815: data = 4'd8;
		11'd816: data = 4'd3;
		11'd817: data = 4'd2;
		11'd818: data = 4'd1;
		11'd819: data = 4'd1;
		11'd820: data = 4'd1;
		11'd821: data = 4'd0;
		11'd822: data = 4'd0;
		11'd823: data = 4'd0;
		11'd824: data = 4'd0;
		11'd825: data = 4'd2;
		11'd826: data = 4'd5;
		11'd827: data = 4'd6;
		11'd828: data = 4'd7;
		11'd829: data = 4'd8;
		11'd830: data = 4'd9;
		11'd831: data = 4'd9;
		11'd832: data = 4'd3;
		11'd833: data = 4'd2;
		11'd834: data = 4'd1;
		11'd835: data = 4'd1;
		11'd836: data = 4'd1;
		11'd837: data = 4'd1;
		11'd838: data = 4'd0;
		11'd839: data = 4'd1;
		11'd840: data = 4'd0;
		11'd841: data = 4'd1;
		11'd842: data = 4'd3;
		11'd843: data = 4'd6;
		11'd844: data = 4'd7;
		11'd845: data = 4'd8;
		11'd846: data = 4'd8;
		11'd847: data = 4'd9;
		11'd848: data = 4'd0;
		11'd849: data = 4'd0;
		11'd850: data = 4'd1;
		11'd851: data = 4'd1;
		11'd852: data = 4'd2;
		11'd853: data = 4'd5;
		11'd854: data = 4'd6;
		11'd855: data = 4'd8;
		11'd856: data = 4'd3;
		11'd857: data = 4'd2;
		11'd858: data = 4'd1;
		11'd859: data = 4'd0;
		11'd860: data = 4'd1;
		11'd861: data = 4'd0;
		11'd862: data = 4'd0;
		11'd863: data = 4'd0;
		11'd864: data = 4'd0;
		11'd865: data = 4'd0;
		11'd866: data = 4'd1;
		11'd867: data = 4'd2;
		11'd868: data = 4'd2;
		11'd869: data = 4'd3;
		11'd870: data = 4'd5;
		11'd871: data = 4'd6;
		11'd872: data = 4'd4;
		11'd873: data = 4'd3;
		11'd874: data = 4'd2;
		11'd875: data = 4'd1;
		11'd876: data = 4'd1;
		11'd877: data = 4'd1;
		11'd878: data = 4'd0;
		11'd879: data = 4'd0;
		11'd880: data = 4'd4;
		11'd881: data = 4'd3;
		11'd882: data = 4'd2;
		11'd883: data = 4'd1;
		11'd884: data = 4'd1;
		11'd885: data = 4'd1;
		11'd886: data = 4'd1;
		11'd887: data = 4'd0;
		11'd888: data = 4'd3;
		11'd889: data = 4'd2;
		11'd890: data = 4'd2;
		11'd891: data = 4'd1;
		11'd892: data = 4'd0;
		11'd893: data = 4'd0;
		11'd894: data = 4'd0;
		11'd895: data = 4'd0;
		11'd896: data = 4'd0;
		11'd897: data = 4'd2;
		11'd898: data = 4'd4;
		11'd899: data = 4'd4;
		11'd900: data = 4'd6;
		11'd901: data = 4'd7;
		11'd902: data = 4'd8;
		11'd903: data = 4'd9;
		11'd904: data = 4'd0;
		11'd905: data = 4'd1;
		11'd906: data = 4'd2;
		11'd907: data = 4'd3;
		11'd908: data = 4'd4;
		11'd909: data = 4'd6;
		11'd910: data = 4'd7;
		11'd911: data = 4'd8;
		11'd912: data = 4'd0;
		11'd913: data = 4'd1;
		11'd914: data = 4'd1;
		11'd915: data = 4'd2;
		11'd916: data = 4'd2;
		11'd917: data = 4'd4;
		11'd918: data = 4'd7;
		11'd919: data = 4'd8;
		11'd920: data = 4'd0;
		11'd921: data = 4'd0;
		11'd922: data = 4'd0;
		11'd923: data = 4'd1;
		11'd924: data = 4'd1;
		11'd925: data = 4'd2;
		11'd926: data = 4'd4;
		11'd927: data = 4'd6;
		11'd928: data = 4'd1;
		11'd929: data = 4'd0;
		11'd930: data = 4'd1;
		11'd931: data = 4'd1;
		11'd932: data = 4'd1;
		11'd933: data = 4'd1;
		11'd934: data = 4'd3;
		11'd935: data = 4'd5;
		11'd936: data = 4'd2;
		11'd937: data = 4'd0;
		11'd938: data = 4'd1;
		11'd939: data = 4'd1;
		11'd940: data = 4'd1;
		11'd941: data = 4'd1;
		11'd942: data = 4'd2;
		11'd943: data = 4'd4;
		11'd944: data = 4'd0;
		11'd945: data = 4'd2;
		11'd946: data = 4'd3;
		11'd947: data = 4'd3;
		11'd948: data = 4'd4;
		11'd949: data = 4'd4;
		11'd950: data = 4'd4;
		11'd951: data = 4'd4;
		11'd952: data = 4'd2;
		11'd953: data = 4'd0;
		11'd954: data = 4'd0;
		11'd955: data = 4'd1;
		11'd956: data = 4'd0;
		11'd957: data = 4'd0;
		11'd958: data = 4'd1;
		11'd959: data = 4'd1;
		11'd960: data = 4'd3;
		11'd961: data = 4'd1;
		11'd962: data = 4'd0;
		11'd963: data = 4'd1;
		11'd964: data = 4'd1;
		11'd965: data = 4'd0;
		11'd966: data = 4'd1;
		11'd967: data = 4'd1;
		11'd968: data = 4'd0;
		11'd969: data = 4'd0;
		11'd970: data = 4'd3;
		11'd971: data = 4'd5;
		11'd972: data = 4'd7;
		11'd973: data = 4'd7;
		11'd974: data = 4'd7;
		11'd975: data = 4'd7;
		11'd976: data = 4'd3;
		11'd977: data = 4'd1;
		11'd978: data = 4'd0;
		11'd979: data = 4'd0;
		11'd980: data = 4'd0;
		11'd981: data = 4'd0;
		11'd982: data = 4'd0;
		11'd983: data = 4'd1;
		11'd984: data = 4'd0;
		11'd985: data = 4'd0;
		11'd986: data = 4'd1;
		11'd987: data = 4'd3;
		11'd988: data = 4'd5;
		11'd989: data = 4'd6;
		11'd990: data = 4'd7;
		11'd991: data = 4'd7;
		11'd992: data = 4'd3;
		11'd993: data = 4'd2;
		11'd994: data = 4'd1;
		11'd995: data = 4'd0;
		11'd996: data = 4'd0;
		11'd997: data = 4'd0;
		11'd998: data = 4'd0;
		11'd999: data = 4'd1;
		11'd1000: data = 4'd0;
		11'd1001: data = 4'd1;
		11'd1002: data = 4'd1;
		11'd1003: data = 4'd2;
		11'd1004: data = 4'd3;
		11'd1005: data = 4'd5;
		11'd1006: data = 4'd6;
		11'd1007: data = 4'd7;
		11'd1008: data = 4'd0;
		11'd1009: data = 4'd1;
		11'd1010: data = 4'd1;
		11'd1011: data = 4'd2;
		11'd1012: data = 4'd3;
		11'd1013: data = 4'd3;
		11'd1014: data = 4'd4;
		11'd1015: data = 4'd6;
		11'd1016: data = 4'd0;
		11'd1017: data = 4'd2;
		11'd1018: data = 4'd4;
		11'd1019: data = 4'd7;
		11'd1020: data = 4'd8;
		11'd1021: data = 4'd8;
		11'd1022: data = 4'd8;
		11'd1023: data = 4'd8;
		11'd1024: data = 4'd0;
		11'd1025: data = 4'd2;
		11'd1026: data = 4'd4;
		11'd1027: data = 4'd7;
		11'd1028: data = 4'd9;
		11'd1029: data = 4'd9;
		11'd1030: data = 4'd9;
		11'd1031: data = 4'd10;
		11'd1032: data = 4'd0;
		11'd1033: data = 4'd1;
		11'd1034: data = 4'd3;
		11'd1035: data = 4'd6;
		11'd1036: data = 4'd8;
		11'd1037: data = 4'd9;
		11'd1038: data = 4'd10;
		11'd1039: data = 4'd10;
		11'd1040: data = 4'd0;
		11'd1041: data = 4'd1;
		11'd1042: data = 4'd2;
		11'd1043: data = 4'd4;
		11'd1044: data = 4'd7;
		11'd1045: data = 4'd9;
		11'd1046: data = 4'd9;
		11'd1047: data = 4'd10;
		11'd1048: data = 4'd0;
		11'd1049: data = 4'd0;
		11'd1050: data = 4'd0;
		11'd1051: data = 4'd1;
		11'd1052: data = 4'd4;
		11'd1053: data = 4'd6;
		11'd1054: data = 4'd8;
		11'd1055: data = 4'd9;
		11'd1056: data = 4'd1;
		11'd1057: data = 4'd0;
		11'd1058: data = 4'd0;
		11'd1059: data = 4'd1;
		11'd1060: data = 4'd2;
		11'd1061: data = 4'd5;
		11'd1062: data = 4'd7;
		11'd1063: data = 4'd9;
		11'd1064: data = 4'd2;
		11'd1065: data = 4'd0;
		11'd1066: data = 4'd1;
		11'd1067: data = 4'd1;
		11'd1068: data = 4'd2;
		11'd1069: data = 4'd3;
		11'd1070: data = 4'd6;
		11'd1071: data = 4'd8;
		11'd1072: data = 4'd2;
		11'd1073: data = 4'd0;
		11'd1074: data = 4'd0;
		11'd1075: data = 4'd0;
		11'd1076: data = 4'd1;
		11'd1077: data = 4'd2;
		11'd1078: data = 4'd2;
		11'd1079: data = 4'd6;
		11'd1080: data = 4'd2;
		11'd1081: data = 4'd1;
		11'd1082: data = 4'd0;
		11'd1083: data = 4'd1;
		11'd1084: data = 4'd1;
		11'd1085: data = 4'd2;
		11'd1086: data = 4'd2;
		11'd1087: data = 4'd3;
		11'd1088: data = 4'd3;
		11'd1089: data = 4'd2;
		11'd1090: data = 4'd0;
		11'd1091: data = 4'd1;
		11'd1092: data = 4'd1;
		11'd1093: data = 4'd1;
		11'd1094: data = 4'd2;
		11'd1095: data = 4'd3;
		11'd1096: data = 4'd0;
		11'd1097: data = 4'd4;
		11'd1098: data = 4'd5;
		11'd1099: data = 4'd6;
		11'd1100: data = 4'd6;
		11'd1101: data = 4'd6;
		11'd1102: data = 4'd6;
		11'd1103: data = 4'd6;
		11'd1104: data = 4'd3;
		11'd1105: data = 4'd2;
		11'd1106: data = 4'd0;
		11'd1107: data = 4'd0;
		11'd1108: data = 4'd0;
		11'd1109: data = 4'd0;
		11'd1110: data = 4'd1;
		11'd1111: data = 4'd2;
		11'd1112: data = 4'd0;
		11'd1113: data = 4'd0;
		11'd1114: data = 4'd3;
		11'd1115: data = 4'd4;
		11'd1116: data = 4'd5;
		11'd1117: data = 4'd5;
		11'd1118: data = 4'd5;
		11'd1119: data = 4'd5;
		11'd1120: data = 4'd3;
		11'd1121: data = 4'd2;
		11'd1122: data = 4'd1;
		11'd1123: data = 4'd0;
		11'd1124: data = 4'd0;
		11'd1125: data = 4'd0;
		11'd1126: data = 4'd1;
		11'd1127: data = 4'd2;
		11'd1128: data = 4'd0;
		11'd1129: data = 4'd1;
		11'd1130: data = 4'd1;
		11'd1131: data = 4'd2;
		11'd1132: data = 4'd2;
		11'd1133: data = 4'd3;
		11'd1134: data = 4'd5;
		11'd1135: data = 4'd5;
		11'd1136: data = 4'd0;
		11'd1137: data = 4'd1;
		11'd1138: data = 4'd2;
		11'd1139: data = 4'd3;
		11'd1140: data = 4'd3;
		11'd1141: data = 4'd4;
		11'd1142: data = 4'd4;
		11'd1143: data = 4'd6;
		11'd1144: data = 4'd5;
		11'd1145: data = 4'd4;
		11'd1146: data = 4'd3;
		11'd1147: data = 4'd2;
		11'd1148: data = 4'd0;
		11'd1149: data = 4'd0;
		11'd1150: data = 4'd1;
		11'd1151: data = 4'd1;
		11'd1152: data = 4'd5;
		11'd1153: data = 4'd4;
		11'd1154: data = 4'd3;
		11'd1155: data = 4'd2;
		11'd1156: data = 4'd1;
		11'd1157: data = 4'd0;
		11'd1158: data = 4'd0;
		11'd1159: data = 4'd1;
		11'd1160: data = 4'd0;
		11'd1161: data = 4'd2;
		11'd1162: data = 4'd6;
		11'd1163: data = 4'd7;
		11'd1164: data = 4'd7;
		11'd1165: data = 4'd7;
		11'd1166: data = 4'd7;
		11'd1167: data = 4'd7;
		11'd1168: data = 4'd0;
		11'd1169: data = 4'd3;
		11'd1170: data = 4'd6;
		11'd1171: data = 4'd10;
		11'd1172: data = 4'd10;
		11'd1173: data = 4'd10;
		11'd1174: data = 4'd10;
		11'd1175: data = 4'd10;
		11'd1176: data = 4'd0;
		11'd1177: data = 4'd1;
		11'd1178: data = 4'd2;
		11'd1179: data = 4'd7;
		11'd1180: data = 4'd11;
		11'd1181: data = 4'd11;
		11'd1182: data = 4'd11;
		11'd1183: data = 4'd11;
		11'd1184: data = 4'd1;
		11'd1185: data = 4'd0;
		11'd1186: data = 4'd1;
		11'd1187: data = 4'd4;
		11'd1188: data = 4'd9;
		11'd1189: data = 4'd11;
		11'd1190: data = 4'd11;
		11'd1191: data = 4'd11;
		11'd1192: data = 4'd1;
		11'd1193: data = 4'd0;
		11'd1194: data = 4'd0;
		11'd1195: data = 4'd1;
		11'd1196: data = 4'd5;
		11'd1197: data = 4'd9;
		11'd1198: data = 4'd10;
		11'd1199: data = 4'd10;
		11'd1200: data = 4'd1;
		11'd1201: data = 4'd0;
		11'd1202: data = 4'd0;
		11'd1203: data = 4'd1;
		11'd1204: data = 4'd3;
		11'd1205: data = 4'd7;
		11'd1206: data = 4'd10;
		11'd1207: data = 4'd10;
		11'd1208: data = 4'd1;
		11'd1209: data = 4'd0;
		11'd1210: data = 4'd0;
		11'd1211: data = 4'd0;
		11'd1212: data = 4'd2;
		11'd1213: data = 4'd3;
		11'd1214: data = 4'd7;
		11'd1215: data = 4'd9;
		11'd1216: data = 4'd2;
		11'd1217: data = 4'd1;
		11'd1218: data = 4'd0;
		11'd1219: data = 4'd0;
		11'd1220: data = 4'd2;
		11'd1221: data = 4'd3;
		11'd1222: data = 4'd4;
		11'd1223: data = 4'd7;
		11'd1224: data = 4'd3;
		11'd1225: data = 4'd2;
		11'd1226: data = 4'd0;
		11'd1227: data = 4'd1;
		11'd1228: data = 4'd2;
		11'd1229: data = 4'd3;
		11'd1230: data = 4'd4;
		11'd1231: data = 4'd4;
		11'd1232: data = 4'd3;
		11'd1233: data = 4'd1;
		11'd1234: data = 4'd0;
		11'd1235: data = 4'd0;
		11'd1236: data = 4'd1;
		11'd1237: data = 4'd2;
		11'd1238: data = 4'd2;
		11'd1239: data = 4'd3;
		11'd1240: data = 4'd0;
		11'd1241: data = 4'd1;
		11'd1242: data = 4'd3;
		11'd1243: data = 4'd4;
		11'd1244: data = 4'd4;
		11'd1245: data = 4'd4;
		11'd1246: data = 4'd4;
		11'd1247: data = 4'd4;
		11'd1248: data = 4'd4;
		11'd1249: data = 4'd3;
		11'd1250: data = 4'd2;
		11'd1251: data = 4'd0;
		11'd1252: data = 4'd0;
		11'd1253: data = 4'd1;
		11'd1254: data = 4'd2;
		11'd1255: data = 4'd3;
		11'd1256: data = 4'd0;
		11'd1257: data = 4'd1;
		11'd1258: data = 4'd1;
		11'd1259: data = 4'd2;
		11'd1260: data = 4'd4;
		11'd1261: data = 4'd4;
		11'd1262: data = 4'd4;
		11'd1263: data = 4'd4;
		11'd1264: data = 4'd5;
		11'd1265: data = 4'd3;
		11'd1266: data = 4'd2;
		11'd1267: data = 4'd1;
		11'd1268: data = 4'd0;
		11'd1269: data = 4'd1;
		11'd1270: data = 4'd2;
		11'd1271: data = 4'd3;
		11'd1272: data = 4'd4;
		11'd1273: data = 4'd3;
		11'd1274: data = 4'd2;
		11'd1275: data = 4'd1;
		11'd1276: data = 4'd0;
		11'd1277: data = 4'd0;
		11'd1278: data = 4'd1;
		11'd1279: data = 4'd1;
		11'd1280: data = 4'd0;
		11'd1281: data = 4'd4;
		11'd1282: data = 4'd8;
		11'd1283: data = 4'd9;
		11'd1284: data = 4'd9;
		11'd1285: data = 4'd9;
		11'd1286: data = 4'd9;
		11'd1287: data = 4'd9;
		11'd1288: data = 4'd0;
		11'd1289: data = 4'd3;
		11'd1290: data = 4'd7;
		11'd1291: data = 4'd11;
		11'd1292: data = 4'd11;
		11'd1293: data = 4'd11;
		11'd1294: data = 4'd11;
		11'd1295: data = 4'd11;
		11'd1296: data = 4'd1;
		11'd1297: data = 4'd0;
		11'd1298: data = 4'd3;
		11'd1299: data = 4'd7;
		11'd1300: data = 4'd11;
		11'd1301: data = 4'd11;
		11'd1302: data = 4'd11;
		11'd1303: data = 4'd11;
		11'd1304: data = 4'd1;
		11'd1305: data = 4'd0;
		11'd1306: data = 4'd1;
		11'd1307: data = 4'd2;
		11'd1308: data = 4'd6;
		11'd1309: data = 4'd10;
		11'd1310: data = 4'd10;
		11'd1311: data = 4'd10;
		11'd1312: data = 4'd1;
		11'd1313: data = 4'd0;
		11'd1314: data = 4'd0;
		11'd1315: data = 4'd1;
		11'd1316: data = 4'd2;
		11'd1317: data = 4'd6;
		11'd1318: data = 4'd9;
		11'd1319: data = 4'd9;
		11'd1320: data = 4'd2;
		11'd1321: data = 4'd1;
		11'd1322: data = 4'd0;
		11'd1323: data = 4'd1;
		11'd1324: data = 4'd2;
		11'd1325: data = 4'd4;
		11'd1326: data = 4'd7;
		11'd1327: data = 4'd9;
		11'd1328: data = 4'd3;
		11'd1329: data = 4'd1;
		11'd1330: data = 4'd0;
		11'd1331: data = 4'd1;
		11'd1332: data = 4'd3;
		11'd1333: data = 4'd4;
		11'd1334: data = 4'd5;
		11'd1335: data = 4'd8;
		11'd1336: data = 4'd3;
		11'd1337: data = 4'd1;
		11'd1338: data = 4'd0;
		11'd1339: data = 4'd0;
		11'd1340: data = 4'd2;
		11'd1341: data = 4'd3;
		11'd1342: data = 4'd4;
		11'd1343: data = 4'd5;
		11'd1344: data = 4'd4;
		11'd1345: data = 4'd2;
		11'd1346: data = 4'd1;
		11'd1347: data = 4'd0;
		11'd1348: data = 4'd2;
		11'd1349: data = 4'd3;
		11'd1350: data = 4'd4;
		11'd1351: data = 4'd4;
		11'd1352: data = 4'd4;
		11'd1353: data = 4'd3;
		11'd1354: data = 4'd1;
		11'd1355: data = 4'd0;
		11'd1356: data = 4'd2;
		11'd1357: data = 4'd2;
		11'd1358: data = 4'd3;
		11'd1359: data = 4'd4;
		11'd1360: data = 4'd4;
		11'd1361: data = 4'd3;
		11'd1362: data = 4'd1;
		11'd1363: data = 4'd0;
		11'd1364: data = 4'd0;
		11'd1365: data = 4'd1;
		11'd1366: data = 4'd2;
		11'd1367: data = 4'd3;
		11'd1368: data = 4'd4;
		11'd1369: data = 4'd3;
		11'd1370: data = 4'd2;
		11'd1371: data = 4'd0;
		11'd1372: data = 4'd0;
		11'd1373: data = 4'd0;
		11'd1374: data = 4'd1;
		11'd1375: data = 4'd2;
		11'd1376: data = 4'd0;
		11'd1377: data = 4'd1;
		11'd1378: data = 4'd1;
		11'd1379: data = 4'd2;
		11'd1380: data = 4'd3;
		11'd1381: data = 4'd3;
		11'd1382: data = 4'd3;
		11'd1383: data = 4'd3;
		11'd1384: data = 4'd0;
		11'd1385: data = 4'd3;
		11'd1386: data = 4'd6;
		11'd1387: data = 4'd6;
		11'd1388: data = 4'd6;
		11'd1389: data = 4'd6;
		11'd1390: data = 4'd6;
		11'd1391: data = 4'd6;
		11'd1392: data = 4'd0;
		11'd1393: data = 4'd4;
		11'd1394: data = 4'd7;
		11'd1395: data = 4'd9;
		11'd1396: data = 4'd9;
		11'd1397: data = 4'd9;
		11'd1398: data = 4'd9;
		11'd1399: data = 4'd9;
		11'd1400: data = 4'd0;
		11'd1401: data = 4'd3;
		11'd1402: data = 4'd7;
		11'd1403: data = 4'd10;
		11'd1404: data = 4'd10;
		11'd1405: data = 4'd10;
		11'd1406: data = 4'd10;
		11'd1407: data = 4'd10;
		11'd1408: data = 4'd0;
		11'd1409: data = 4'd1;
		11'd1410: data = 4'd5;
		11'd1411: data = 4'd8;
		11'd1412: data = 4'd10;
		11'd1413: data = 4'd10;
		11'd1414: data = 4'd10;
		11'd1415: data = 4'd10;
		11'd1416: data = 4'd0;
		11'd1417: data = 4'd0;
		11'd1418: data = 4'd3;
		11'd1419: data = 4'd7;
		11'd1420: data = 4'd10;
		11'd1421: data = 4'd10;
		11'd1422: data = 4'd10;
		11'd1423: data = 4'd10;
		11'd1424: data = 4'd1;
		11'd1425: data = 4'd0;
		11'd1426: data = 4'd1;
		11'd1427: data = 4'd4;
		11'd1428: data = 4'd8;
		11'd1429: data = 4'd10;
		11'd1430: data = 4'd10;
		11'd1431: data = 4'd10;
		11'd1432: data = 4'd1;
		11'd1433: data = 4'd0;
		11'd1434: data = 4'd0;
		11'd1435: data = 4'd2;
		11'd1436: data = 4'd5;
		11'd1437: data = 4'd9;
		11'd1438: data = 4'd9;
		11'd1439: data = 4'd9;
		11'd1440: data = 4'd1;
		11'd1441: data = 4'd0;
		11'd1442: data = 4'd0;
		11'd1443: data = 4'd1;
		11'd1444: data = 4'd2;
		11'd1445: data = 4'd4;
		11'd1446: data = 4'd8;
		11'd1447: data = 4'd8;
		11'd1448: data = 4'd2;
		11'd1449: data = 4'd0;
		11'd1450: data = 4'd0;
		11'd1451: data = 4'd1;
		11'd1452: data = 4'd2;
		11'd1453: data = 4'd4;
		11'd1454: data = 4'd5;
		11'd1455: data = 4'd8;
		11'd1456: data = 4'd2;
		11'd1457: data = 4'd1;
		11'd1458: data = 4'd0;
		11'd1459: data = 4'd1;
		11'd1460: data = 4'd2;
		11'd1461: data = 4'd4;
		11'd1462: data = 4'd5;
		11'd1463: data = 4'd6;
		11'd1464: data = 4'd2;
		11'd1465: data = 4'd1;
		11'd1466: data = 4'd0;
		11'd1467: data = 4'd0;
		11'd1468: data = 4'd1;
		11'd1469: data = 4'd3;
		11'd1470: data = 4'd4;
		11'd1471: data = 4'd5;
		11'd1472: data = 4'd0;
		11'd1473: data = 4'd2;
		11'd1474: data = 4'd2;
		11'd1475: data = 4'd2;
		11'd1476: data = 4'd2;
		11'd1477: data = 4'd2;
		11'd1478: data = 4'd2;
		11'd1479: data = 4'd2;
		11'd1480: data = 4'd3;
		11'd1481: data = 4'd2;
		11'd1482: data = 4'd0;
		11'd1483: data = 4'd0;
		11'd1484: data = 4'd1;
		11'd1485: data = 4'd3;
		11'd1486: data = 4'd4;
		11'd1487: data = 4'd4;
		11'd1488: data = 4'd3;
		11'd1489: data = 4'd2;
		11'd1490: data = 4'd0;
		11'd1491: data = 4'd0;
		11'd1492: data = 4'd1;
		11'd1493: data = 4'd2;
		11'd1494: data = 4'd2;
		11'd1495: data = 4'd3;
		default: data = 4'd0;
	endcase
end
endmodule

module layer0_N24_idx_1(address, data);
input wire [8:0] address;
output reg [7:0] data;

always @(*) begin
	case(address)
		9'd0: data = 8'd0;
		9'd1: data = 8'd0;
		9'd2: data = 8'd0;
		9'd3: data = 8'd0;
		9'd4: data = 8'd0;
		9'd5: data = 8'd0;
		9'd6: data = 8'd0;
		9'd7: data = 8'd0;
		9'd8: data = 8'd0;
		9'd9: data = 8'd0;
		9'd10: data = 8'd0;
		9'd11: data = 8'd0;
		9'd12: data = 8'd0;
		9'd13: data = 8'd0;
		9'd14: data = 8'd0;
		9'd15: data = 8'd0;
		9'd16: data = 8'd0;
		9'd17: data = 8'd0;
		9'd18: data = 8'd0;
		9'd19: data = 8'd0;
		9'd20: data = 8'd0;
		9'd21: data = 8'd0;
		9'd22: data = 8'd0;
		9'd23: data = 8'd0;
		9'd24: data = 8'd0;
		9'd25: data = 8'd0;
		9'd26: data = 8'd0;
		9'd27: data = 8'd0;
		9'd28: data = 8'd0;
		9'd29: data = 8'd0;
		9'd30: data = 8'd0;
		9'd31: data = 8'd0;
		9'd32: data = 8'd0;
		9'd33: data = 8'd0;
		9'd34: data = 8'd0;
		9'd35: data = 8'd0;
		9'd36: data = 8'd0;
		9'd37: data = 8'd0;
		9'd38: data = 8'd0;
		9'd39: data = 8'd0;
		9'd40: data = 8'd0;
		9'd41: data = 8'd0;
		9'd42: data = 8'd0;
		9'd43: data = 8'd0;
		9'd44: data = 8'd0;
		9'd45: data = 8'd0;
		9'd46: data = 8'd0;
		9'd47: data = 8'd0;
		9'd48: data = 8'd0;
		9'd49: data = 8'd0;
		9'd50: data = 8'd0;
		9'd51: data = 8'd0;
		9'd52: data = 8'd0;
		9'd53: data = 8'd0;
		9'd54: data = 8'd0;
		9'd55: data = 8'd0;
		9'd56: data = 8'd0;
		9'd57: data = 8'd0;
		9'd58: data = 8'd0;
		9'd59: data = 8'd0;
		9'd60: data = 8'd0;
		9'd61: data = 8'd0;
		9'd62: data = 8'd0;
		9'd63: data = 8'd0;
		9'd64: data = 8'd0;
		9'd65: data = 8'd9;
		9'd66: data = 8'd0;
		9'd67: data = 8'd9;
		9'd68: data = 8'd0;
		9'd69: data = 8'd0;
		9'd70: data = 8'd0;
		9'd71: data = 8'd0;
		9'd72: data = 8'd0;
		9'd73: data = 8'd0;
		9'd74: data = 8'd0;
		9'd75: data = 8'd0;
		9'd76: data = 8'd0;
		9'd77: data = 8'd0;
		9'd78: data = 8'd0;
		9'd79: data = 8'd0;
		9'd80: data = 8'd0;
		9'd81: data = 8'd0;
		9'd82: data = 8'd0;
		9'd83: data = 8'd0;
		9'd84: data = 8'd0;
		9'd85: data = 8'd0;
		9'd86: data = 8'd0;
		9'd87: data = 8'd0;
		9'd88: data = 8'd0;
		9'd89: data = 8'd0;
		9'd90: data = 8'd0;
		9'd91: data = 8'd0;
		9'd92: data = 8'd0;
		9'd93: data = 8'd0;
		9'd94: data = 8'd0;
		9'd95: data = 8'd0;
		9'd96: data = 8'd0;
		9'd97: data = 8'd10;
		9'd98: data = 8'd0;
		9'd99: data = 8'd44;
		9'd100: data = 8'd0;
		9'd101: data = 8'd10;
		9'd102: data = 8'd0;
		9'd103: data = 8'd26;
		9'd104: data = 8'd0;
		9'd105: data = 8'd0;
		9'd106: data = 8'd0;
		9'd107: data = 8'd9;
		9'd108: data = 8'd0;
		9'd109: data = 8'd0;
		9'd110: data = 8'd0;
		9'd111: data = 8'd0;
		9'd112: data = 8'd0;
		9'd113: data = 8'd0;
		9'd114: data = 8'd0;
		9'd115: data = 8'd0;
		9'd116: data = 8'd0;
		9'd117: data = 8'd0;
		9'd118: data = 8'd0;
		9'd119: data = 8'd0;
		9'd120: data = 8'd0;
		9'd121: data = 8'd9;
		9'd122: data = 8'd0;
		9'd123: data = 8'd9;
		9'd124: data = 8'd0;
		9'd125: data = 8'd0;
		9'd126: data = 8'd0;
		9'd127: data = 8'd0;
		9'd128: data = 8'd0;
		9'd129: data = 8'd27;
		9'd130: data = 8'd0;
		9'd131: data = 8'd16;
		9'd132: data = 8'd0;
		9'd133: data = 8'd45;
		9'd134: data = 8'd0;
		9'd135: data = 8'd17;
		9'd136: data = 8'd0;
		9'd137: data = 8'd0;
		9'd138: data = 8'd0;
		9'd139: data = 8'd16;
		9'd140: data = 8'd0;
		9'd141: data = 8'd10;
		9'd142: data = 8'd0;
		9'd143: data = 8'd4;
		9'd144: data = 8'd0;
		9'd145: data = 8'd4;
		9'd146: data = 8'd0;
		9'd147: data = 8'd4;
		9'd148: data = 8'd0;
		9'd149: data = 8'd4;
		9'd150: data = 8'd0;
		9'd151: data = 8'd4;
		9'd152: data = 8'd0;
		9'd153: data = 8'd10;
		9'd154: data = 8'd0;
		9'd155: data = 8'd10;
		9'd156: data = 8'd0;
		9'd157: data = 8'd26;
		9'd158: data = 8'd0;
		9'd159: data = 8'd0;
		9'd160: data = 8'd0;
		9'd161: data = 8'd18;
		9'd162: data = 8'd0;
		9'd163: data = 8'd12;
		9'd164: data = 8'd0;
		9'd165: data = 8'd7;
		9'd166: data = 8'd0;
		9'd167: data = 8'd46;
		9'd168: data = 8'd0;
		9'd169: data = 8'd4;
		9'd170: data = 8'd0;
		9'd171: data = 8'd28;
		9'd172: data = 8'd0;
		9'd173: data = 8'd27;
		9'd174: data = 8'd0;
		9'd175: data = 8'd7;
		9'd176: data = 8'd0;
		9'd177: data = 8'd7;
		9'd178: data = 8'd0;
		9'd179: data = 8'd7;
		9'd180: data = 8'd0;
		9'd181: data = 8'd7;
		9'd182: data = 8'd0;
		9'd183: data = 8'd7;
		9'd184: data = 8'd0;
		9'd185: data = 8'd17;
		9'd186: data = 8'd0;
		9'd187: data = 8'd17;
		9'd188: data = 8'd0;
		9'd189: data = 8'd0;
		9'd190: data = 8'd0;
		9'd191: data = 8'd16;
		9'd192: data = 8'd0;
		9'd193: data = 8'd19;
		9'd194: data = 8'd0;
		9'd195: data = 8'd47;
		9'd196: data = 8'd0;
		9'd197: data = 8'd48;
		9'd198: data = 8'd0;
		9'd199: data = 8'd29;
		9'd200: data = 8'd0;
		9'd201: data = 8'd49;
		9'd202: data = 8'd0;
		9'd203: data = 8'd50;
		9'd204: data = 8'd0;
		9'd205: data = 8'd51;
		9'd206: data = 8'd0;
		9'd207: data = 8'd13;
		9'd208: data = 8'd0;
		9'd209: data = 8'd13;
		9'd210: data = 8'd0;
		9'd211: data = 8'd18;
		9'd212: data = 8'd0;
		9'd213: data = 8'd18;
		9'd214: data = 8'd0;
		9'd215: data = 8'd13;
		9'd216: data = 8'd0;
		9'd217: data = 8'd13;
		9'd218: data = 8'd1;
		9'd219: data = 8'd12;
		9'd220: data = 8'd1;
		9'd221: data = 8'd12;
		9'd222: data = 8'd5;
		9'd223: data = 8'd28;
		9'd224: data = 8'd0;
		9'd225: data = 8'd30;
		9'd226: data = 8'd0;
		9'd227: data = 8'd11;
		9'd228: data = 8'd0;
		9'd229: data = 8'd20;
		9'd230: data = 8'd0;
		9'd231: data = 8'd31;
		9'd232: data = 8'd0;
		9'd233: data = 8'd52;
		9'd234: data = 8'd0;
		9'd235: data = 8'd53;
		9'd236: data = 8'd0;
		9'd237: data = 8'd29;
		9'd238: data = 8'd1;
		9'd239: data = 8'd54;
		9'd240: data = 8'd1;
		9'd241: data = 8'd55;
		9'd242: data = 8'd5;
		9'd243: data = 8'd8;
		9'd244: data = 8'd5;
		9'd245: data = 8'd8;
		9'd246: data = 8'd3;
		9'd247: data = 8'd32;
		9'd248: data = 8'd3;
		9'd249: data = 8'd8;
		9'd250: data = 8'd1;
		9'd251: data = 8'd8;
		9'd252: data = 8'd1;
		9'd253: data = 8'd56;
		9'd254: data = 8'd57;
		9'd255: data = 8'd58;
		9'd256: data = 8'd59;
		9'd257: data = 8'd33;
		9'd258: data = 8'd4;
		9'd259: data = 8'd33;
		9'd260: data = 8'd12;
		9'd261: data = 8'd34;
		9'd262: data = 8'd60;
		9'd263: data = 8'd61;
		9'd264: data = 8'd62;
		9'd265: data = 8'd20;
		9'd266: data = 8'd63;
		9'd267: data = 8'd64;
		9'd268: data = 8'd65;
		9'd269: data = 8'd66;
		9'd270: data = 8'd21;
		9'd271: data = 8'd67;
		9'd272: data = 8'd68;
		9'd273: data = 8'd69;
		9'd274: data = 8'd5;
		9'd275: data = 8'd70;
		9'd276: data = 8'd3;
		9'd277: data = 8'd8;
		9'd278: data = 8'd3;
		9'd279: data = 8'd8;
		9'd280: data = 8'd1;
		9'd281: data = 8'd32;
		9'd282: data = 8'd1;
		9'd283: data = 8'd71;
		9'd284: data = 8'd22;
		9'd285: data = 8'd19;
		9'd286: data = 8'd22;
		9'd287: data = 8'd19;
		9'd288: data = 8'd72;
		9'd289: data = 8'd35;
		9'd290: data = 8'd73;
		9'd291: data = 8'd74;
		9'd292: data = 8'd75;
		9'd293: data = 8'd35;
		9'd294: data = 8'd0;
		9'd295: data = 8'd76;
		9'd296: data = 8'd77;
		9'd297: data = 8'd78;
		9'd298: data = 8'd79;
		9'd299: data = 8'd80;
		9'd300: data = 8'd21;
		9'd301: data = 8'd81;
		9'd302: data = 8'd82;
		9'd303: data = 8'd83;
		9'd304: data = 8'd84;
		9'd305: data = 8'd36;
		9'd306: data = 8'd85;
		9'd307: data = 8'd86;
		9'd308: data = 8'd87;
		9'd309: data = 8'd88;
		9'd310: data = 8'd5;
		9'd311: data = 8'd89;
		9'd312: data = 8'd3;
		9'd313: data = 8'd11;
		9'd314: data = 8'd3;
		9'd315: data = 8'd11;
		9'd316: data = 8'd90;
		9'd317: data = 8'd11;
		9'd318: data = 8'd1;
		9'd319: data = 8'd11;
		9'd320: data = 8'd91;
		9'd321: data = 8'd14;
		9'd322: data = 8'd92;
		9'd323: data = 8'd93;
		9'd324: data = 8'd94;
		9'd325: data = 8'd95;
		9'd326: data = 8'd96;
		9'd327: data = 8'd97;
		9'd328: data = 8'd98;
		9'd329: data = 8'd23;
		9'd330: data = 8'd99;
		9'd331: data = 8'd100;
		9'd332: data = 8'd21;
		9'd333: data = 8'd101;
		9'd334: data = 8'd102;
		9'd335: data = 8'd103;
		9'd336: data = 8'd104;
		9'd337: data = 8'd105;
		9'd338: data = 8'd5;
		9'd339: data = 8'd36;
		9'd340: data = 8'd3;
		9'd341: data = 8'd106;
		9'd342: data = 8'd107;
		9'd343: data = 8'd108;
		9'd344: data = 8'd109;
		9'd345: data = 8'd20;
		9'd346: data = 8'd110;
		9'd347: data = 8'd37;
		9'd348: data = 8'd111;
		9'd349: data = 8'd37;
		9'd350: data = 8'd1;
		9'd351: data = 8'd30;
		9'd352: data = 8'd14;
		9'd353: data = 8'd2;
		9'd354: data = 8'd112;
		9'd355: data = 8'd6;
		9'd356: data = 8'd113;
		9'd357: data = 8'd38;
		9'd358: data = 8'd114;
		9'd359: data = 8'd25;
		9'd360: data = 8'd115;
		9'd361: data = 8'd15;
		9'd362: data = 8'd116;
		9'd363: data = 8'd15;
		9'd364: data = 8'd117;
		9'd365: data = 8'd118;
		9'd366: data = 8'd119;
		9'd367: data = 8'd38;
		9'd368: data = 8'd120;
		9'd369: data = 8'd15;
		9'd370: data = 8'd5;
		9'd371: data = 8'd121;
		9'd372: data = 8'd122;
		9'd373: data = 8'd123;
		9'd374: data = 8'd124;
		9'd375: data = 8'd125;
		9'd376: data = 8'd3;
		9'd377: data = 8'd126;
		9'd378: data = 8'd1;
		9'd379: data = 8'd39;
		9'd380: data = 8'd1;
		9'd381: data = 8'd39;
		9'd382: data = 8'd22;
		9'd383: data = 8'd40;
		9'd384: data = 8'd127;
		9'd385: data = 8'd0;
		9'd386: data = 8'd128;
		9'd387: data = 8'd0;
		9'd388: data = 8'd129;
		9'd389: data = 8'd0;
		9'd390: data = 8'd130;
		9'd391: data = 8'd0;
		9'd392: data = 8'd131;
		9'd393: data = 8'd2;
		9'd394: data = 8'd132;
		9'd395: data = 8'd2;
		9'd396: data = 8'd133;
		9'd397: data = 8'd2;
		9'd398: data = 8'd134;
		9'd399: data = 8'd2;
		9'd400: data = 8'd135;
		9'd401: data = 8'd2;
		9'd402: data = 8'd136;
		9'd403: data = 8'd137;
		9'd404: data = 8'd138;
		9'd405: data = 8'd139;
		9'd406: data = 8'd140;
		9'd407: data = 8'd42;
		9'd408: data = 8'd24;
		9'd409: data = 8'd141;
		9'd410: data = 8'd24;
		9'd411: data = 8'd142;
		9'd412: data = 8'd143;
		9'd413: data = 8'd40;
		9'd414: data = 8'd144;
		9'd415: data = 8'd23;
		9'd416: data = 8'd145;
		9'd417: data = 8'd0;
		9'd418: data = 8'd146;
		9'd419: data = 8'd0;
		9'd420: data = 8'd25;
		9'd421: data = 8'd0;
		9'd422: data = 8'd147;
		9'd423: data = 8'd0;
		9'd424: data = 8'd148;
		9'd425: data = 8'd0;
		9'd426: data = 8'd149;
		9'd427: data = 8'd0;
		9'd428: data = 8'd150;
		9'd429: data = 8'd0;
		9'd430: data = 8'd151;
		9'd431: data = 8'd0;
		9'd432: data = 8'd152;
		9'd433: data = 8'd0;
		9'd434: data = 8'd153;
		9'd435: data = 8'd2;
		9'd436: data = 8'd154;
		9'd437: data = 8'd6;
		9'd438: data = 8'd41;
		9'd439: data = 8'd155;
		9'd440: data = 8'd156;
		9'd441: data = 8'd157;
		9'd442: data = 8'd158;
		9'd443: data = 8'd34;
		9'd444: data = 8'd24;
		9'd445: data = 8'd31;
		9'd446: data = 8'd159;
		9'd447: data = 8'd23;
		9'd448: data = 8'd2;
		9'd449: data = 8'd0;
		9'd450: data = 8'd160;
		9'd451: data = 8'd0;
		9'd452: data = 8'd161;
		9'd453: data = 8'd0;
		9'd454: data = 8'd25;
		9'd455: data = 8'd0;
		9'd456: data = 8'd162;
		9'd457: data = 8'd0;
		9'd458: data = 8'd42;
		9'd459: data = 8'd0;
		9'd460: data = 8'd163;
		9'd461: data = 8'd0;
		9'd462: data = 8'd164;
		9'd463: data = 8'd0;
		9'd464: data = 8'd165;
		9'd465: data = 8'd0;
		9'd466: data = 8'd166;
		9'd467: data = 8'd0;
		9'd468: data = 8'd167;
		9'd469: data = 8'd2;
		9'd470: data = 8'd168;
		9'd471: data = 8'd2;
		9'd472: data = 8'd169;
		9'd473: data = 8'd15;
		9'd474: data = 8'd170;
		9'd475: data = 8'd14;
		9'd476: data = 8'd43;
		9'd477: data = 8'd14;
		9'd478: data = 8'd171;
		9'd479: data = 8'd172;
		9'd480: data = 8'd6;
		9'd481: data = 8'd0;
		9'd482: data = 8'd173;
		9'd483: data = 8'd0;
		9'd484: data = 8'd174;
		9'd485: data = 8'd0;
		9'd486: data = 8'd175;
		9'd487: data = 8'd0;
		9'd488: data = 8'd176;
		9'd489: data = 8'd0;
		9'd490: data = 8'd177;
		9'd491: data = 8'd0;
		9'd492: data = 8'd178;
		9'd493: data = 8'd0;
		9'd494: data = 8'd179;
		9'd495: data = 8'd0;
		9'd496: data = 8'd180;
		9'd497: data = 8'd0;
		9'd498: data = 8'd181;
		9'd499: data = 8'd0;
		9'd500: data = 8'd182;
		9'd501: data = 8'd0;
		9'd502: data = 8'd183;
		9'd503: data = 8'd184;
		9'd504: data = 8'd185;
		9'd505: data = 8'd6;
		9'd506: data = 8'd186;
		9'd507: data = 8'd6;
		9'd508: data = 8'd41;
		9'd509: data = 8'd6;
		9'd510: data = 8'd43;
		9'd511: data = 8'd6;
		default: data = 8'd0;
	endcase
end
endmodule

module layer0_N24_rsh_1(address, data);
input wire [8:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		9'd0: data = 2'd3;
		9'd1: data = 2'd3;
		9'd2: data = 2'd3;
		9'd3: data = 2'd3;
		9'd4: data = 2'd3;
		9'd5: data = 2'd3;
		9'd6: data = 2'd3;
		9'd7: data = 2'd3;
		9'd8: data = 2'd3;
		9'd9: data = 2'd3;
		9'd10: data = 2'd3;
		9'd11: data = 2'd3;
		9'd12: data = 2'd3;
		9'd13: data = 2'd3;
		9'd14: data = 2'd3;
		9'd15: data = 2'd3;
		9'd16: data = 2'd3;
		9'd17: data = 2'd3;
		9'd18: data = 2'd3;
		9'd19: data = 2'd3;
		9'd20: data = 2'd3;
		9'd21: data = 2'd3;
		9'd22: data = 2'd3;
		9'd23: data = 2'd3;
		9'd24: data = 2'd3;
		9'd25: data = 2'd3;
		9'd26: data = 2'd3;
		9'd27: data = 2'd3;
		9'd28: data = 2'd3;
		9'd29: data = 2'd3;
		9'd30: data = 2'd3;
		9'd31: data = 2'd3;
		9'd32: data = 2'd3;
		9'd33: data = 2'd2;
		9'd34: data = 2'd3;
		9'd35: data = 2'd3;
		9'd36: data = 2'd3;
		9'd37: data = 2'd3;
		9'd38: data = 2'd3;
		9'd39: data = 2'd3;
		9'd40: data = 2'd3;
		9'd41: data = 2'd3;
		9'd42: data = 2'd3;
		9'd43: data = 2'd3;
		9'd44: data = 2'd3;
		9'd45: data = 2'd3;
		9'd46: data = 2'd3;
		9'd47: data = 2'd3;
		9'd48: data = 2'd3;
		9'd49: data = 2'd3;
		9'd50: data = 2'd3;
		9'd51: data = 2'd3;
		9'd52: data = 2'd3;
		9'd53: data = 2'd3;
		9'd54: data = 2'd3;
		9'd55: data = 2'd3;
		9'd56: data = 2'd3;
		9'd57: data = 2'd3;
		9'd58: data = 2'd3;
		9'd59: data = 2'd3;
		9'd60: data = 2'd3;
		9'd61: data = 2'd3;
		9'd62: data = 2'd3;
		9'd63: data = 2'd3;
		9'd64: data = 2'd3;
		9'd65: data = 2'd0;
		9'd66: data = 2'd3;
		9'd67: data = 2'd1;
		9'd68: data = 2'd3;
		9'd69: data = 2'd2;
		9'd70: data = 2'd3;
		9'd71: data = 2'd2;
		9'd72: data = 2'd3;
		9'd73: data = 2'd2;
		9'd74: data = 2'd3;
		9'd75: data = 2'd3;
		9'd76: data = 2'd3;
		9'd77: data = 2'd3;
		9'd78: data = 2'd3;
		9'd79: data = 2'd3;
		9'd80: data = 2'd3;
		9'd81: data = 2'd3;
		9'd82: data = 2'd3;
		9'd83: data = 2'd3;
		9'd84: data = 2'd3;
		9'd85: data = 2'd2;
		9'd86: data = 2'd3;
		9'd87: data = 2'd3;
		9'd88: data = 2'd3;
		9'd89: data = 2'd3;
		9'd90: data = 2'd3;
		9'd91: data = 2'd3;
		9'd92: data = 2'd3;
		9'd93: data = 2'd3;
		9'd94: data = 2'd3;
		9'd95: data = 2'd3;
		9'd96: data = 2'd3;
		9'd97: data = 2'd0;
		9'd98: data = 2'd3;
		9'd99: data = 2'd0;
		9'd100: data = 2'd3;
		9'd101: data = 2'd1;
		9'd102: data = 2'd3;
		9'd103: data = 2'd0;
		9'd104: data = 2'd3;
		9'd105: data = 2'd1;
		9'd106: data = 2'd3;
		9'd107: data = 2'd1;
		9'd108: data = 2'd3;
		9'd109: data = 2'd2;
		9'd110: data = 2'd3;
		9'd111: data = 2'd2;
		9'd112: data = 2'd3;
		9'd113: data = 2'd1;
		9'd114: data = 2'd3;
		9'd115: data = 2'd1;
		9'd116: data = 2'd3;
		9'd117: data = 2'd1;
		9'd118: data = 2'd3;
		9'd119: data = 2'd1;
		9'd120: data = 2'd3;
		9'd121: data = 2'd1;
		9'd122: data = 2'd3;
		9'd123: data = 2'd1;
		9'd124: data = 2'd3;
		9'd125: data = 2'd2;
		9'd126: data = 2'd3;
		9'd127: data = 2'd2;
		9'd128: data = 2'd3;
		9'd129: data = 2'd0;
		9'd130: data = 2'd3;
		9'd131: data = 2'd0;
		9'd132: data = 2'd3;
		9'd133: data = 2'd0;
		9'd134: data = 2'd3;
		9'd135: data = 2'd0;
		9'd136: data = 2'd3;
		9'd137: data = 2'd0;
		9'd138: data = 2'd3;
		9'd139: data = 2'd1;
		9'd140: data = 2'd3;
		9'd141: data = 2'd1;
		9'd142: data = 2'd3;
		9'd143: data = 2'd1;
		9'd144: data = 2'd3;
		9'd145: data = 2'd1;
		9'd146: data = 2'd3;
		9'd147: data = 2'd1;
		9'd148: data = 2'd3;
		9'd149: data = 2'd1;
		9'd150: data = 2'd3;
		9'd151: data = 2'd1;
		9'd152: data = 2'd3;
		9'd153: data = 2'd1;
		9'd154: data = 2'd3;
		9'd155: data = 2'd1;
		9'd156: data = 2'd3;
		9'd157: data = 2'd0;
		9'd158: data = 2'd3;
		9'd159: data = 2'd1;
		9'd160: data = 2'd3;
		9'd161: data = 2'd0;
		9'd162: data = 2'd3;
		9'd163: data = 2'd0;
		9'd164: data = 2'd3;
		9'd165: data = 2'd0;
		9'd166: data = 2'd3;
		9'd167: data = 2'd0;
		9'd168: data = 2'd3;
		9'd169: data = 2'd0;
		9'd170: data = 2'd3;
		9'd171: data = 2'd0;
		9'd172: data = 2'd3;
		9'd173: data = 2'd1;
		9'd174: data = 2'd3;
		9'd175: data = 2'd1;
		9'd176: data = 2'd3;
		9'd177: data = 2'd1;
		9'd178: data = 2'd3;
		9'd179: data = 2'd1;
		9'd180: data = 2'd3;
		9'd181: data = 2'd1;
		9'd182: data = 2'd3;
		9'd183: data = 2'd1;
		9'd184: data = 2'd3;
		9'd185: data = 2'd0;
		9'd186: data = 2'd3;
		9'd187: data = 2'd0;
		9'd188: data = 2'd3;
		9'd189: data = 2'd0;
		9'd190: data = 2'd3;
		9'd191: data = 2'd1;
		9'd192: data = 2'd3;
		9'd193: data = 2'd0;
		9'd194: data = 2'd3;
		9'd195: data = 2'd0;
		9'd196: data = 2'd3;
		9'd197: data = 2'd0;
		9'd198: data = 2'd3;
		9'd199: data = 2'd0;
		9'd200: data = 2'd3;
		9'd201: data = 2'd0;
		9'd202: data = 2'd3;
		9'd203: data = 2'd0;
		9'd204: data = 2'd3;
		9'd205: data = 2'd0;
		9'd206: data = 2'd3;
		9'd207: data = 2'd0;
		9'd208: data = 2'd3;
		9'd209: data = 2'd0;
		9'd210: data = 2'd3;
		9'd211: data = 2'd1;
		9'd212: data = 2'd3;
		9'd213: data = 2'd1;
		9'd214: data = 2'd3;
		9'd215: data = 2'd0;
		9'd216: data = 2'd3;
		9'd217: data = 2'd0;
		9'd218: data = 2'd2;
		9'd219: data = 2'd1;
		9'd220: data = 2'd2;
		9'd221: data = 2'd1;
		9'd222: data = 2'd0;
		9'd223: data = 2'd0;
		9'd224: data = 2'd2;
		9'd225: data = 2'd0;
		9'd226: data = 2'd3;
		9'd227: data = 2'd0;
		9'd228: data = 2'd3;
		9'd229: data = 2'd0;
		9'd230: data = 2'd3;
		9'd231: data = 2'd0;
		9'd232: data = 2'd3;
		9'd233: data = 2'd0;
		9'd234: data = 2'd3;
		9'd235: data = 2'd0;
		9'd236: data = 2'd3;
		9'd237: data = 2'd0;
		9'd238: data = 2'd2;
		9'd239: data = 2'd0;
		9'd240: data = 2'd2;
		9'd241: data = 2'd0;
		9'd242: data = 2'd0;
		9'd243: data = 2'd0;
		9'd244: data = 2'd0;
		9'd245: data = 2'd0;
		9'd246: data = 2'd0;
		9'd247: data = 2'd0;
		9'd248: data = 2'd0;
		9'd249: data = 2'd0;
		9'd250: data = 2'd0;
		9'd251: data = 2'd0;
		9'd252: data = 2'd0;
		9'd253: data = 2'd0;
		9'd254: data = 2'd0;
		9'd255: data = 2'd0;
		9'd256: data = 2'd0;
		9'd257: data = 2'd0;
		9'd258: data = 2'd1;
		9'd259: data = 2'd0;
		9'd260: data = 2'd2;
		9'd261: data = 2'd0;
		9'd262: data = 2'd0;
		9'd263: data = 2'd0;
		9'd264: data = 2'd0;
		9'd265: data = 2'd0;
		9'd266: data = 2'd0;
		9'd267: data = 2'd0;
		9'd268: data = 2'd0;
		9'd269: data = 2'd0;
		9'd270: data = 2'd0;
		9'd271: data = 2'd0;
		9'd272: data = 2'd0;
		9'd273: data = 2'd0;
		9'd274: data = 2'd0;
		9'd275: data = 2'd0;
		9'd276: data = 2'd0;
		9'd277: data = 2'd0;
		9'd278: data = 2'd0;
		9'd279: data = 2'd0;
		9'd280: data = 2'd0;
		9'd281: data = 2'd0;
		9'd282: data = 2'd0;
		9'd283: data = 2'd0;
		9'd284: data = 2'd0;
		9'd285: data = 2'd1;
		9'd286: data = 2'd0;
		9'd287: data = 2'd1;
		9'd288: data = 2'd0;
		9'd289: data = 2'd0;
		9'd290: data = 2'd0;
		9'd291: data = 2'd0;
		9'd292: data = 2'd0;
		9'd293: data = 2'd0;
		9'd294: data = 2'd1;
		9'd295: data = 2'd0;
		9'd296: data = 2'd0;
		9'd297: data = 2'd0;
		9'd298: data = 2'd0;
		9'd299: data = 2'd0;
		9'd300: data = 2'd0;
		9'd301: data = 2'd0;
		9'd302: data = 2'd0;
		9'd303: data = 2'd0;
		9'd304: data = 2'd0;
		9'd305: data = 2'd0;
		9'd306: data = 2'd0;
		9'd307: data = 2'd0;
		9'd308: data = 2'd0;
		9'd309: data = 2'd0;
		9'd310: data = 2'd0;
		9'd311: data = 2'd0;
		9'd312: data = 2'd0;
		9'd313: data = 2'd1;
		9'd314: data = 2'd0;
		9'd315: data = 2'd1;
		9'd316: data = 2'd0;
		9'd317: data = 2'd1;
		9'd318: data = 2'd0;
		9'd319: data = 2'd1;
		9'd320: data = 2'd0;
		9'd321: data = 2'd1;
		9'd322: data = 2'd0;
		9'd323: data = 2'd0;
		9'd324: data = 2'd0;
		9'd325: data = 2'd0;
		9'd326: data = 2'd0;
		9'd327: data = 2'd0;
		9'd328: data = 2'd0;
		9'd329: data = 2'd0;
		9'd330: data = 2'd0;
		9'd331: data = 2'd0;
		9'd332: data = 2'd0;
		9'd333: data = 2'd0;
		9'd334: data = 2'd0;
		9'd335: data = 2'd0;
		9'd336: data = 2'd0;
		9'd337: data = 2'd0;
		9'd338: data = 2'd0;
		9'd339: data = 2'd0;
		9'd340: data = 2'd0;
		9'd341: data = 2'd0;
		9'd342: data = 2'd0;
		9'd343: data = 2'd0;
		9'd344: data = 2'd0;
		9'd345: data = 2'd1;
		9'd346: data = 2'd0;
		9'd347: data = 2'd0;
		9'd348: data = 2'd0;
		9'd349: data = 2'd0;
		9'd350: data = 2'd0;
		9'd351: data = 2'd1;
		9'd352: data = 2'd0;
		9'd353: data = 2'd2;
		9'd354: data = 2'd0;
		9'd355: data = 2'd1;
		9'd356: data = 2'd0;
		9'd357: data = 2'd1;
		9'd358: data = 2'd0;
		9'd359: data = 2'd2;
		9'd360: data = 2'd0;
		9'd361: data = 2'd1;
		9'd362: data = 2'd0;
		9'd363: data = 2'd1;
		9'd364: data = 2'd0;
		9'd365: data = 2'd0;
		9'd366: data = 2'd0;
		9'd367: data = 2'd0;
		9'd368: data = 2'd0;
		9'd369: data = 2'd0;
		9'd370: data = 2'd0;
		9'd371: data = 2'd0;
		9'd372: data = 2'd0;
		9'd373: data = 2'd0;
		9'd374: data = 2'd0;
		9'd375: data = 2'd0;
		9'd376: data = 2'd0;
		9'd377: data = 2'd0;
		9'd378: data = 2'd0;
		9'd379: data = 2'd0;
		9'd380: data = 2'd0;
		9'd381: data = 2'd0;
		9'd382: data = 2'd0;
		9'd383: data = 2'd0;
		9'd384: data = 2'd0;
		9'd385: data = 2'd3;
		9'd386: data = 2'd0;
		9'd387: data = 2'd3;
		9'd388: data = 2'd0;
		9'd389: data = 2'd3;
		9'd390: data = 2'd0;
		9'd391: data = 2'd3;
		9'd392: data = 2'd0;
		9'd393: data = 2'd2;
		9'd394: data = 2'd0;
		9'd395: data = 2'd2;
		9'd396: data = 2'd0;
		9'd397: data = 2'd2;
		9'd398: data = 2'd0;
		9'd399: data = 2'd2;
		9'd400: data = 2'd0;
		9'd401: data = 2'd1;
		9'd402: data = 2'd0;
		9'd403: data = 2'd0;
		9'd404: data = 2'd0;
		9'd405: data = 2'd0;
		9'd406: data = 2'd0;
		9'd407: data = 2'd1;
		9'd408: data = 2'd0;
		9'd409: data = 2'd0;
		9'd410: data = 2'd0;
		9'd411: data = 2'd0;
		9'd412: data = 2'd0;
		9'd413: data = 2'd0;
		9'd414: data = 2'd0;
		9'd415: data = 2'd0;
		9'd416: data = 2'd0;
		9'd417: data = 2'd3;
		9'd418: data = 2'd0;
		9'd419: data = 2'd3;
		9'd420: data = 2'd0;
		9'd421: data = 2'd3;
		9'd422: data = 2'd0;
		9'd423: data = 2'd3;
		9'd424: data = 2'd0;
		9'd425: data = 2'd3;
		9'd426: data = 2'd0;
		9'd427: data = 2'd3;
		9'd428: data = 2'd0;
		9'd429: data = 2'd3;
		9'd430: data = 2'd0;
		9'd431: data = 2'd3;
		9'd432: data = 2'd0;
		9'd433: data = 2'd3;
		9'd434: data = 2'd0;
		9'd435: data = 2'd2;
		9'd436: data = 2'd0;
		9'd437: data = 2'd0;
		9'd438: data = 2'd0;
		9'd439: data = 2'd0;
		9'd440: data = 2'd0;
		9'd441: data = 2'd0;
		9'd442: data = 2'd0;
		9'd443: data = 2'd1;
		9'd444: data = 2'd0;
		9'd445: data = 2'd1;
		9'd446: data = 2'd0;
		9'd447: data = 2'd0;
		9'd448: data = 2'd0;
		9'd449: data = 2'd3;
		9'd450: data = 2'd0;
		9'd451: data = 2'd3;
		9'd452: data = 2'd0;
		9'd453: data = 2'd3;
		9'd454: data = 2'd0;
		9'd455: data = 2'd3;
		9'd456: data = 2'd0;
		9'd457: data = 2'd3;
		9'd458: data = 2'd0;
		9'd459: data = 2'd3;
		9'd460: data = 2'd0;
		9'd461: data = 2'd3;
		9'd462: data = 2'd0;
		9'd463: data = 2'd3;
		9'd464: data = 2'd0;
		9'd465: data = 2'd3;
		9'd466: data = 2'd0;
		9'd467: data = 2'd3;
		9'd468: data = 2'd0;
		9'd469: data = 2'd2;
		9'd470: data = 2'd0;
		9'd471: data = 2'd1;
		9'd472: data = 2'd0;
		9'd473: data = 2'd1;
		9'd474: data = 2'd0;
		9'd475: data = 2'd1;
		9'd476: data = 2'd0;
		9'd477: data = 2'd1;
		9'd478: data = 2'd0;
		9'd479: data = 2'd0;
		9'd480: data = 2'd0;
		9'd481: data = 2'd3;
		9'd482: data = 2'd0;
		9'd483: data = 2'd3;
		9'd484: data = 2'd0;
		9'd485: data = 2'd3;
		9'd486: data = 2'd0;
		9'd487: data = 2'd3;
		9'd488: data = 2'd0;
		9'd489: data = 2'd3;
		9'd490: data = 2'd0;
		9'd491: data = 2'd3;
		9'd492: data = 2'd0;
		9'd493: data = 2'd3;
		9'd494: data = 2'd0;
		9'd495: data = 2'd3;
		9'd496: data = 2'd0;
		9'd497: data = 2'd3;
		9'd498: data = 2'd0;
		9'd499: data = 2'd3;
		9'd500: data = 2'd0;
		9'd501: data = 2'd3;
		9'd502: data = 2'd0;
		9'd503: data = 2'd0;
		9'd504: data = 2'd0;
		9'd505: data = 2'd1;
		9'd506: data = 2'd0;
		9'd507: data = 2'd1;
		9'd508: data = 2'd0;
		9'd509: data = 2'd1;
		9'd510: data = 2'd0;
		9'd511: data = 2'd1;
		default: data = 2'd0;
	endcase
end
endmodule

module layer0_N24(address, data);
input wire [11:0] address;
output reg [3:0] data;

wire [7:0] i; layer0_N24_idx_1 idx_1_inst(address[11:3], i);
wire [1:0] t; layer0_N24_rsh_1 rsh_1_inst(address[11:3], t);
wire [3:0] b; layer0_N24_2 layer0_N24_2_inst(address[11:3], b);
wire [3:0] u; layer0_N24_ust_1 ust_1_inst({i, address[2:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule
