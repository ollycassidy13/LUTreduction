
module layer1_N3_bias_4(address, data);
input wire [0:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		1'd0: data = 2'd3;
		1'd1: data = 2'd2;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N3_4(address, data);
input wire [3:0] address;
output reg [1:0] data;

wire [1:0] b; layer1_N3_bias_4 bias_4_inst(address[3:3], b);


always @(*) begin
	data = b;
end
endmodule

module layer1_N3_ust_3(address, data);
input wire [3:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		4'd0: data = 3'd0;
		4'd1: data = 3'd3;
		4'd2: data = 3'd3;
		4'd3: data = 3'd6;
		4'd4: data = 3'd0;
		4'd5: data = 3'd2;
		4'd6: data = 3'd2;
		4'd7: data = 3'd3;
		4'd8: data = 3'd0;
		4'd9: data = 3'd2;
		4'd10: data = 3'd2;
		4'd11: data = 3'd4;
		4'd12: data = 3'd0;
		4'd13: data = 3'd3;
		4'd14: data = 3'd3;
		4'd15: data = 3'd5;
		default: data = 3'd0;
	endcase
end
endmodule

module layer1_N3_idx_3(address, data);
input wire [3:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		4'd0: data = 2'd1;
		4'd1: data = 2'd1;
		4'd2: data = 2'd1;
		4'd3: data = 2'd1;
		4'd4: data = 2'd2;
		4'd5: data = 2'd2;
		4'd6: data = 2'd2;
		4'd7: data = 2'd2;
		4'd8: data = 2'd3;
		4'd9: data = 2'd3;
		4'd10: data = 2'd3;
		4'd11: data = 2'd0;
		4'd12: data = 2'd0;
		4'd13: data = 2'd0;
		4'd14: data = 2'd0;
		4'd15: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N3_3(address, data);
input wire [5:0] address;
output reg [3:0] data;

wire [1:0] i; layer1_N3_idx_3 idx_3_inst(address[5:2], i);
wire [1:0] b; layer1_N3_4 layer1_N3_4_inst(address[5:2], b);
wire [2:0] u; layer1_N3_ust_3 ust_3_inst({i, address[1:0]}, u);

always @(*) begin
	data = u + b;
end
endmodule

module layer1_N3_ust_2(address, data);
input wire [7:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		8'd0: data = 3'd0;
		8'd1: data = 3'd0;
		8'd2: data = 3'd0;
		8'd3: data = 3'd0;
		8'd4: data = 3'd0;
		8'd5: data = 3'd1;
		8'd6: data = 3'd1;
		8'd7: data = 3'd2;
		8'd8: data = 3'd0;
		8'd9: data = 3'd0;
		8'd10: data = 3'd0;
		8'd11: data = 3'd1;
		8'd12: data = 3'd1;
		8'd13: data = 3'd2;
		8'd14: data = 3'd2;
		8'd15: data = 3'd3;
		8'd16: data = 3'd0;
		8'd17: data = 3'd1;
		8'd18: data = 3'd0;
		8'd19: data = 3'd1;
		8'd20: data = 3'd0;
		8'd21: data = 3'd1;
		8'd22: data = 3'd0;
		8'd23: data = 3'd0;
		8'd24: data = 3'd0;
		8'd25: data = 3'd0;
		8'd26: data = 3'd1;
		8'd27: data = 3'd2;
		8'd28: data = 3'd2;
		8'd29: data = 3'd3;
		8'd30: data = 3'd3;
		8'd31: data = 3'd4;
		8'd32: data = 3'd0;
		8'd33: data = 3'd2;
		8'd34: data = 3'd0;
		8'd35: data = 3'd2;
		8'd36: data = 3'd1;
		8'd37: data = 3'd3;
		8'd38: data = 3'd1;
		8'd39: data = 3'd3;
		8'd40: data = 3'd0;
		8'd41: data = 3'd1;
		8'd42: data = 3'd1;
		8'd43: data = 3'd2;
		8'd44: data = 3'd2;
		8'd45: data = 3'd3;
		8'd46: data = 3'd3;
		8'd47: data = 3'd4;
		8'd48: data = 3'd0;
		8'd49: data = 3'd1;
		8'd50: data = 3'd0;
		8'd51: data = 3'd1;
		8'd52: data = 3'd0;
		8'd53: data = 3'd0;
		8'd54: data = 3'd0;
		8'd55: data = 3'd0;
		8'd56: data = 3'd0;
		8'd57: data = 3'd0;
		8'd58: data = 3'd1;
		8'd59: data = 3'd1;
		8'd60: data = 3'd1;
		8'd61: data = 3'd2;
		8'd62: data = 3'd2;
		8'd63: data = 3'd3;
		8'd64: data = 3'd0;
		8'd65: data = 3'd2;
		8'd66: data = 3'd1;
		8'd67: data = 3'd3;
		8'd68: data = 3'd1;
		8'd69: data = 3'd3;
		8'd70: data = 3'd2;
		8'd71: data = 3'd4;
		8'd72: data = 3'd1;
		8'd73: data = 3'd1;
		8'd74: data = 3'd0;
		8'd75: data = 3'd1;
		8'd76: data = 3'd0;
		8'd77: data = 3'd1;
		8'd78: data = 3'd0;
		8'd79: data = 3'd1;
		8'd80: data = 3'd0;
		8'd81: data = 3'd1;
		8'd82: data = 3'd0;
		8'd83: data = 3'd2;
		8'd84: data = 3'd1;
		8'd85: data = 3'd3;
		8'd86: data = 3'd2;
		8'd87: data = 3'd4;
		8'd88: data = 3'd0;
		8'd89: data = 3'd1;
		8'd90: data = 3'd1;
		8'd91: data = 3'd2;
		8'd92: data = 3'd1;
		8'd93: data = 3'd3;
		8'd94: data = 3'd2;
		8'd95: data = 3'd4;
		8'd96: data = 3'd0;
		8'd97: data = 3'd0;
		8'd98: data = 3'd0;
		8'd99: data = 3'd0;
		8'd100: data = 3'd1;
		8'd101: data = 3'd2;
		8'd102: data = 3'd2;
		8'd103: data = 3'd3;
		8'd104: data = 3'd0;
		8'd105: data = 3'd1;
		8'd106: data = 3'd1;
		8'd107: data = 3'd2;
		8'd108: data = 3'd2;
		8'd109: data = 3'd4;
		8'd110: data = 3'd3;
		8'd111: data = 3'd5;
		8'd112: data = 3'd0;
		8'd113: data = 3'd1;
		8'd114: data = 3'd1;
		8'd115: data = 3'd1;
		8'd116: data = 3'd0;
		8'd117: data = 3'd1;
		8'd118: data = 3'd0;
		8'd119: data = 3'd1;
		8'd120: data = 3'd0;
		8'd121: data = 3'd0;
		8'd122: data = 3'd0;
		8'd123: data = 3'd0;
		8'd124: data = 3'd0;
		8'd125: data = 3'd1;
		8'd126: data = 3'd0;
		8'd127: data = 3'd2;
		8'd128: data = 3'd0;
		8'd129: data = 3'd2;
		8'd130: data = 3'd1;
		8'd131: data = 3'd2;
		8'd132: data = 3'd1;
		8'd133: data = 3'd3;
		8'd134: data = 3'd2;
		8'd135: data = 3'd4;
		8'd136: data = 3'd0;
		8'd137: data = 3'd1;
		8'd138: data = 3'd0;
		8'd139: data = 3'd2;
		8'd140: data = 3'd1;
		8'd141: data = 3'd3;
		8'd142: data = 3'd1;
		8'd143: data = 3'd3;
		8'd144: data = 3'd0;
		8'd145: data = 3'd1;
		8'd146: data = 3'd1;
		8'd147: data = 3'd3;
		8'd148: data = 3'd2;
		8'd149: data = 3'd4;
		8'd150: data = 3'd2;
		8'd151: data = 3'd4;
		8'd152: data = 3'd0;
		8'd153: data = 3'd1;
		8'd154: data = 3'd1;
		8'd155: data = 3'd3;
		8'd156: data = 3'd2;
		8'd157: data = 3'd4;
		8'd158: data = 3'd3;
		8'd159: data = 3'd5;
		8'd160: data = 3'd0;
		8'd161: data = 3'd2;
		8'd162: data = 3'd1;
		8'd163: data = 3'd3;
		8'd164: data = 3'd2;
		8'd165: data = 3'd4;
		8'd166: data = 3'd3;
		8'd167: data = 3'd5;
		8'd168: data = 3'd0;
		8'd169: data = 3'd0;
		8'd170: data = 3'd0;
		8'd171: data = 3'd0;
		8'd172: data = 3'd0;
		8'd173: data = 3'd1;
		8'd174: data = 3'd1;
		8'd175: data = 3'd3;
		8'd176: data = 3'd0;
		8'd177: data = 3'd1;
		8'd178: data = 3'd1;
		8'd179: data = 3'd2;
		8'd180: data = 3'd2;
		8'd181: data = 3'd3;
		8'd182: data = 3'd2;
		8'd183: data = 3'd4;
		8'd184: data = 3'd0;
		8'd185: data = 3'd1;
		8'd186: data = 3'd1;
		8'd187: data = 3'd2;
		8'd188: data = 3'd2;
		8'd189: data = 3'd3;
		8'd190: data = 3'd3;
		8'd191: data = 3'd5;
		default: data = 3'd0;
	endcase
end
endmodule

module layer1_N3_idx_2(address, data);
input wire [5:0] address;
output reg [4:0] data;

always @(*) begin
	case(address)
		6'd0: data = 5'd7;
		6'd1: data = 5'd14;
		6'd2: data = 5'd15;
		6'd3: data = 5'd4;
		6'd4: data = 5'd7;
		6'd5: data = 5'd4;
		6'd6: data = 5'd0;
		6'd7: data = 5'd16;
		6'd8: data = 5'd1;
		6'd9: data = 5'd4;
		6'd10: data = 5'd0;
		6'd11: data = 5'd8;
		6'd12: data = 5'd1;
		6'd13: data = 5'd9;
		6'd14: data = 5'd0;
		6'd15: data = 5'd8;
		6'd16: data = 5'd1;
		6'd17: data = 5'd9;
		6'd18: data = 5'd0;
		6'd19: data = 5'd17;
		6'd20: data = 5'd1;
		6'd21: data = 5'd4;
		6'd22: data = 5'd0;
		6'd23: data = 5'd10;
		6'd24: data = 5'd1;
		6'd25: data = 5'd2;
		6'd26: data = 5'd0;
		6'd27: data = 5'd10;
		6'd28: data = 5'd1;
		6'd29: data = 5'd2;
		6'd30: data = 5'd0;
		6'd31: data = 5'd11;
		6'd32: data = 5'd5;
		6'd33: data = 5'd2;
		6'd34: data = 5'd0;
		6'd35: data = 5'd18;
		6'd36: data = 5'd5;
		6'd37: data = 5'd2;
		6'd38: data = 5'd0;
		6'd39: data = 5'd19;
		6'd40: data = 5'd5;
		6'd41: data = 5'd2;
		6'd42: data = 5'd0;
		6'd43: data = 5'd20;
		6'd44: data = 5'd3;
		6'd45: data = 5'd2;
		6'd46: data = 5'd0;
		6'd47: data = 5'd11;
		6'd48: data = 5'd3;
		6'd49: data = 5'd2;
		6'd50: data = 5'd21;
		6'd51: data = 5'd22;
		6'd52: data = 5'd3;
		6'd53: data = 5'd6;
		6'd54: data = 5'd12;
		6'd55: data = 5'd23;
		6'd56: data = 5'd3;
		6'd57: data = 5'd6;
		6'd58: data = 5'd12;
		6'd59: data = 5'd13;
		6'd60: data = 5'd3;
		6'd61: data = 5'd6;
		6'd62: data = 5'd1;
		6'd63: data = 5'd13;
		default: data = 5'd0;
	endcase
end
endmodule

module layer1_N3_rsh_2(address, data);
input wire [5:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		6'd0: data = 1'd0;
		6'd1: data = 1'd0;
		6'd2: data = 1'd0;
		6'd3: data = 1'd0;
		6'd4: data = 1'd0;
		6'd5: data = 1'd1;
		6'd6: data = 1'd0;
		6'd7: data = 1'd0;
		6'd8: data = 1'd0;
		6'd9: data = 1'd1;
		6'd10: data = 1'd0;
		6'd11: data = 1'd0;
		6'd12: data = 1'd0;
		6'd13: data = 1'd0;
		6'd14: data = 1'd0;
		6'd15: data = 1'd0;
		6'd16: data = 1'd0;
		6'd17: data = 1'd0;
		6'd18: data = 1'd0;
		6'd19: data = 1'd0;
		6'd20: data = 1'd0;
		6'd21: data = 1'd1;
		6'd22: data = 1'd0;
		6'd23: data = 1'd0;
		6'd24: data = 1'd0;
		6'd25: data = 1'd0;
		6'd26: data = 1'd0;
		6'd27: data = 1'd0;
		6'd28: data = 1'd0;
		6'd29: data = 1'd0;
		6'd30: data = 1'd0;
		6'd31: data = 1'd0;
		6'd32: data = 1'd0;
		6'd33: data = 1'd0;
		6'd34: data = 1'd0;
		6'd35: data = 1'd0;
		6'd36: data = 1'd0;
		6'd37: data = 1'd0;
		6'd38: data = 1'd0;
		6'd39: data = 1'd0;
		6'd40: data = 1'd0;
		6'd41: data = 1'd0;
		6'd42: data = 1'd0;
		6'd43: data = 1'd0;
		6'd44: data = 1'd0;
		6'd45: data = 1'd0;
		6'd46: data = 1'd0;
		6'd47: data = 1'd0;
		6'd48: data = 1'd0;
		6'd49: data = 1'd0;
		6'd50: data = 1'd0;
		6'd51: data = 1'd0;
		6'd52: data = 1'd0;
		6'd53: data = 1'd0;
		6'd54: data = 1'd0;
		6'd55: data = 1'd0;
		6'd56: data = 1'd0;
		6'd57: data = 1'd0;
		6'd58: data = 1'd0;
		6'd59: data = 1'd0;
		6'd60: data = 1'd0;
		6'd61: data = 1'd0;
		6'd62: data = 1'd0;
		6'd63: data = 1'd0;
		default: data = 1'd0;
	endcase
end
endmodule

module layer1_N3_2(address, data);
input wire [8:0] address;
output reg [3:0] data;

wire [4:0] i; layer1_N3_idx_2 idx_2_inst(address[8:3], i);
wire [0:0] t; layer1_N3_rsh_2 rsh_2_inst(address[8:3], t);
wire [3:0] b; layer1_N3_3 layer1_N3_3_inst(address[8:3], b);
wire [2:0] u; layer1_N3_ust_2 ust_2_inst({i, address[2:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule

module layer1_N3_ust_1(address, data);
input wire [7:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		8'd0: data = 2'd0;
		8'd1: data = 2'd0;
		8'd2: data = 2'd0;
		8'd3: data = 2'd0;
		8'd4: data = 2'd1;
		8'd5: data = 2'd1;
		8'd6: data = 2'd1;
		8'd7: data = 2'd1;
		8'd8: data = 2'd0;
		8'd9: data = 2'd1;
		8'd10: data = 2'd1;
		8'd11: data = 2'd1;
		8'd12: data = 2'd1;
		8'd13: data = 2'd2;
		8'd14: data = 2'd2;
		8'd15: data = 2'd2;
		8'd16: data = 2'd0;
		8'd17: data = 2'd0;
		8'd18: data = 2'd0;
		8'd19: data = 2'd1;
		8'd20: data = 2'd1;
		8'd21: data = 2'd1;
		8'd22: data = 2'd1;
		8'd23: data = 2'd1;
		8'd24: data = 2'd0;
		8'd25: data = 2'd0;
		8'd26: data = 2'd1;
		8'd27: data = 2'd1;
		8'd28: data = 2'd1;
		8'd29: data = 2'd1;
		8'd30: data = 2'd2;
		8'd31: data = 2'd2;
		8'd32: data = 2'd0;
		8'd33: data = 2'd0;
		8'd34: data = 2'd1;
		8'd35: data = 2'd1;
		8'd36: data = 2'd1;
		8'd37: data = 2'd1;
		8'd38: data = 2'd1;
		8'd39: data = 2'd1;
		8'd40: data = 2'd0;
		8'd41: data = 2'd0;
		8'd42: data = 2'd0;
		8'd43: data = 2'd1;
		8'd44: data = 2'd1;
		8'd45: data = 2'd1;
		8'd46: data = 2'd1;
		8'd47: data = 2'd2;
		8'd48: data = 2'd0;
		8'd49: data = 2'd1;
		8'd50: data = 2'd1;
		8'd51: data = 2'd1;
		8'd52: data = 2'd1;
		8'd53: data = 2'd1;
		8'd54: data = 2'd1;
		8'd55: data = 2'd1;
		8'd56: data = 2'd0;
		8'd57: data = 2'd1;
		8'd58: data = 2'd1;
		8'd59: data = 2'd1;
		8'd60: data = 2'd1;
		8'd61: data = 2'd1;
		8'd62: data = 2'd2;
		8'd63: data = 2'd2;
		8'd64: data = 2'd0;
		8'd65: data = 2'd0;
		8'd66: data = 2'd0;
		8'd67: data = 2'd0;
		8'd68: data = 2'd0;
		8'd69: data = 2'd1;
		8'd70: data = 2'd1;
		8'd71: data = 2'd0;
		8'd72: data = 2'd0;
		8'd73: data = 2'd1;
		8'd74: data = 2'd1;
		8'd75: data = 2'd1;
		8'd76: data = 2'd1;
		8'd77: data = 2'd1;
		8'd78: data = 2'd1;
		8'd79: data = 2'd2;
		8'd80: data = 2'd0;
		8'd81: data = 2'd0;
		8'd82: data = 2'd1;
		8'd83: data = 2'd1;
		8'd84: data = 2'd1;
		8'd85: data = 2'd1;
		8'd86: data = 2'd1;
		8'd87: data = 2'd2;
		8'd88: data = 2'd1;
		8'd89: data = 2'd0;
		8'd90: data = 2'd0;
		8'd91: data = 2'd0;
		8'd92: data = 2'd0;
		8'd93: data = 2'd0;
		8'd94: data = 2'd0;
		8'd95: data = 2'd0;
		8'd96: data = 2'd1;
		8'd97: data = 2'd1;
		8'd98: data = 2'd1;
		8'd99: data = 2'd0;
		8'd100: data = 2'd0;
		8'd101: data = 2'd0;
		8'd102: data = 2'd0;
		8'd103: data = 2'd0;
		8'd104: data = 2'd1;
		8'd105: data = 2'd1;
		8'd106: data = 2'd0;
		8'd107: data = 2'd0;
		8'd108: data = 2'd0;
		8'd109: data = 2'd0;
		8'd110: data = 2'd0;
		8'd111: data = 2'd0;
		8'd112: data = 2'd0;
		8'd113: data = 2'd0;
		8'd114: data = 2'd0;
		8'd115: data = 2'd0;
		8'd116: data = 2'd0;
		8'd117: data = 2'd0;
		8'd118: data = 2'd1;
		8'd119: data = 2'd0;
		8'd120: data = 2'd1;
		8'd121: data = 2'd0;
		8'd122: data = 2'd1;
		8'd123: data = 2'd1;
		8'd124: data = 2'd1;
		8'd125: data = 2'd1;
		8'd126: data = 2'd1;
		8'd127: data = 2'd1;
		8'd128: data = 2'd1;
		8'd129: data = 2'd1;
		8'd130: data = 2'd1;
		8'd131: data = 2'd1;
		8'd132: data = 2'd1;
		8'd133: data = 2'd1;
		8'd134: data = 2'd0;
		8'd135: data = 2'd1;
		8'd136: data = 2'd1;
		8'd137: data = 2'd1;
		8'd138: data = 2'd1;
		8'd139: data = 2'd1;
		8'd140: data = 2'd0;
		8'd141: data = 2'd0;
		8'd142: data = 2'd0;
		8'd143: data = 2'd1;
		8'd144: data = 2'd1;
		8'd145: data = 2'd1;
		8'd146: data = 2'd1;
		8'd147: data = 2'd0;
		8'd148: data = 2'd0;
		8'd149: data = 2'd0;
		8'd150: data = 2'd0;
		8'd151: data = 2'd1;
		8'd152: data = 2'd1;
		8'd153: data = 2'd1;
		8'd154: data = 2'd0;
		8'd155: data = 2'd0;
		8'd156: data = 2'd0;
		8'd157: data = 2'd0;
		8'd158: data = 2'd0;
		8'd159: data = 2'd1;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N3_idx_1(address, data);
input wire [8:0] address;
output reg [4:0] data;

always @(*) begin
	case(address)
		9'd0: data = 5'd0;
		9'd1: data = 5'd12;
		9'd2: data = 5'd0;
		9'd3: data = 5'd0;
		9'd4: data = 5'd0;
		9'd5: data = 5'd0;
		9'd6: data = 5'd3;
		9'd7: data = 5'd0;
		9'd8: data = 5'd6;
		9'd9: data = 5'd0;
		9'd10: data = 5'd0;
		9'd11: data = 5'd0;
		9'd12: data = 5'd4;
		9'd13: data = 5'd0;
		9'd14: data = 5'd0;
		9'd15: data = 5'd0;
		9'd16: data = 5'd8;
		9'd17: data = 5'd4;
		9'd18: data = 5'd0;
		9'd19: data = 5'd0;
		9'd20: data = 5'd5;
		9'd21: data = 5'd0;
		9'd22: data = 5'd9;
		9'd23: data = 5'd0;
		9'd24: data = 5'd2;
		9'd25: data = 5'd0;
		9'd26: data = 5'd1;
		9'd27: data = 5'd4;
		9'd28: data = 5'd2;
		9'd29: data = 5'd0;
		9'd30: data = 5'd1;
		9'd31: data = 5'd3;
		9'd32: data = 5'd0;
		9'd33: data = 5'd13;
		9'd34: data = 5'd0;
		9'd35: data = 5'd0;
		9'd36: data = 5'd0;
		9'd37: data = 5'd0;
		9'd38: data = 5'd3;
		9'd39: data = 5'd0;
		9'd40: data = 5'd6;
		9'd41: data = 5'd0;
		9'd42: data = 5'd6;
		9'd43: data = 5'd0;
		9'd44: data = 5'd4;
		9'd45: data = 5'd0;
		9'd46: data = 5'd0;
		9'd47: data = 5'd0;
		9'd48: data = 5'd14;
		9'd49: data = 5'd2;
		9'd50: data = 5'd0;
		9'd51: data = 5'd0;
		9'd52: data = 5'd5;
		9'd53: data = 5'd0;
		9'd54: data = 5'd3;
		9'd55: data = 5'd0;
		9'd56: data = 5'd5;
		9'd57: data = 5'd0;
		9'd58: data = 5'd1;
		9'd59: data = 5'd6;
		9'd60: data = 5'd10;
		9'd61: data = 5'd2;
		9'd62: data = 5'd0;
		9'd63: data = 5'd0;
		9'd64: data = 5'd1;
		9'd65: data = 5'd11;
		9'd66: data = 5'd15;
		9'd67: data = 5'd0;
		9'd68: data = 5'd1;
		9'd69: data = 5'd0;
		9'd70: data = 5'd1;
		9'd71: data = 5'd0;
		9'd72: data = 5'd6;
		9'd73: data = 5'd0;
		9'd74: data = 5'd6;
		9'd75: data = 5'd0;
		9'd76: data = 5'd2;
		9'd77: data = 5'd0;
		9'd78: data = 5'd1;
		9'd79: data = 5'd0;
		9'd80: data = 5'd0;
		9'd81: data = 5'd1;
		9'd82: data = 5'd0;
		9'd83: data = 5'd0;
		9'd84: data = 5'd3;
		9'd85: data = 5'd0;
		9'd86: data = 5'd3;
		9'd87: data = 5'd0;
		9'd88: data = 5'd3;
		9'd89: data = 5'd0;
		9'd90: data = 5'd0;
		9'd91: data = 5'd5;
		9'd92: data = 5'd3;
		9'd93: data = 5'd4;
		9'd94: data = 5'd5;
		9'd95: data = 5'd2;
		9'd96: data = 5'd1;
		9'd97: data = 5'd0;
		9'd98: data = 5'd2;
		9'd99: data = 5'd0;
		9'd100: data = 5'd1;
		9'd101: data = 5'd0;
		9'd102: data = 5'd1;
		9'd103: data = 5'd0;
		9'd104: data = 5'd0;
		9'd105: data = 5'd0;
		9'd106: data = 5'd4;
		9'd107: data = 5'd0;
		9'd108: data = 5'd2;
		9'd109: data = 5'd0;
		9'd110: data = 5'd1;
		9'd111: data = 5'd0;
		9'd112: data = 5'd0;
		9'd113: data = 5'd3;
		9'd114: data = 5'd0;
		9'd115: data = 5'd0;
		9'd116: data = 5'd3;
		9'd117: data = 5'd0;
		9'd118: data = 5'd3;
		9'd119: data = 5'd0;
		9'd120: data = 5'd7;
		9'd121: data = 5'd0;
		9'd122: data = 5'd2;
		9'd123: data = 5'd3;
		9'd124: data = 5'd1;
		9'd125: data = 5'd7;
		9'd126: data = 5'd3;
		9'd127: data = 5'd10;
		9'd128: data = 5'd8;
		9'd129: data = 5'd0;
		9'd130: data = 5'd2;
		9'd131: data = 5'd0;
		9'd132: data = 5'd0;
		9'd133: data = 5'd0;
		9'd134: data = 5'd0;
		9'd135: data = 5'd0;
		9'd136: data = 5'd0;
		9'd137: data = 5'd0;
		9'd138: data = 5'd4;
		9'd139: data = 5'd0;
		9'd140: data = 5'd0;
		9'd141: data = 5'd0;
		9'd142: data = 5'd3;
		9'd143: data = 5'd0;
		9'd144: data = 5'd0;
		9'd145: data = 5'd5;
		9'd146: data = 5'd0;
		9'd147: data = 5'd0;
		9'd148: data = 5'd3;
		9'd149: data = 5'd0;
		9'd150: data = 5'd1;
		9'd151: data = 5'd0;
		9'd152: data = 5'd1;
		9'd153: data = 5'd0;
		9'd154: data = 5'd5;
		9'd155: data = 5'd1;
		9'd156: data = 5'd0;
		9'd157: data = 5'd0;
		9'd158: data = 5'd1;
		9'd159: data = 5'd7;
		9'd160: data = 5'd8;
		9'd161: data = 5'd0;
		9'd162: data = 5'd2;
		9'd163: data = 5'd0;
		9'd164: data = 5'd0;
		9'd165: data = 5'd0;
		9'd166: data = 5'd0;
		9'd167: data = 5'd0;
		9'd168: data = 5'd6;
		9'd169: data = 5'd0;
		9'd170: data = 5'd2;
		9'd171: data = 5'd0;
		9'd172: data = 5'd1;
		9'd173: data = 5'd0;
		9'd174: data = 5'd5;
		9'd175: data = 5'd0;
		9'd176: data = 5'd0;
		9'd177: data = 5'd0;
		9'd178: data = 5'd0;
		9'd179: data = 5'd0;
		9'd180: data = 5'd1;
		9'd181: data = 5'd0;
		9'd182: data = 5'd1;
		9'd183: data = 5'd0;
		9'd184: data = 5'd1;
		9'd185: data = 5'd5;
		9'd186: data = 5'd3;
		9'd187: data = 5'd2;
		9'd188: data = 5'd5;
		9'd189: data = 5'd2;
		9'd190: data = 5'd0;
		9'd191: data = 5'd0;
		9'd192: data = 5'd0;
		9'd193: data = 5'd0;
		9'd194: data = 5'd2;
		9'd195: data = 5'd0;
		9'd196: data = 5'd0;
		9'd197: data = 5'd0;
		9'd198: data = 5'd2;
		9'd199: data = 5'd0;
		9'd200: data = 5'd6;
		9'd201: data = 5'd0;
		9'd202: data = 5'd2;
		9'd203: data = 5'd0;
		9'd204: data = 5'd1;
		9'd205: data = 5'd0;
		9'd206: data = 5'd0;
		9'd207: data = 5'd6;
		9'd208: data = 5'd0;
		9'd209: data = 5'd0;
		9'd210: data = 5'd0;
		9'd211: data = 5'd0;
		9'd212: data = 5'd1;
		9'd213: data = 5'd0;
		9'd214: data = 5'd1;
		9'd215: data = 5'd0;
		9'd216: data = 5'd1;
		9'd217: data = 5'd3;
		9'd218: data = 5'd1;
		9'd219: data = 5'd4;
		9'd220: data = 5'd3;
		9'd221: data = 5'd4;
		9'd222: data = 5'd5;
		9'd223: data = 5'd2;
		9'd224: data = 5'd0;
		9'd225: data = 5'd0;
		9'd226: data = 5'd0;
		9'd227: data = 5'd0;
		9'd228: data = 5'd0;
		9'd229: data = 5'd0;
		9'd230: data = 5'd2;
		9'd231: data = 5'd0;
		9'd232: data = 5'd4;
		9'd233: data = 5'd0;
		9'd234: data = 5'd0;
		9'd235: data = 5'd0;
		9'd236: data = 5'd3;
		9'd237: data = 5'd0;
		9'd238: data = 5'd0;
		9'd239: data = 5'd4;
		9'd240: data = 5'd0;
		9'd241: data = 5'd0;
		9'd242: data = 5'd0;
		9'd243: data = 5'd0;
		9'd244: data = 5'd1;
		9'd245: data = 5'd0;
		9'd246: data = 5'd0;
		9'd247: data = 5'd5;
		9'd248: data = 5'd0;
		9'd249: data = 5'd0;
		9'd250: data = 5'd0;
		9'd251: data = 5'd6;
		9'd252: data = 5'd1;
		9'd253: data = 5'd6;
		9'd254: data = 5'd3;
		9'd255: data = 5'd4;
		9'd256: data = 5'd6;
		9'd257: data = 5'd0;
		9'd258: data = 5'd0;
		9'd259: data = 5'd0;
		9'd260: data = 5'd0;
		9'd261: data = 5'd0;
		9'd262: data = 5'd2;
		9'd263: data = 5'd0;
		9'd264: data = 5'd2;
		9'd265: data = 5'd0;
		9'd266: data = 5'd0;
		9'd267: data = 5'd0;
		9'd268: data = 5'd3;
		9'd269: data = 5'd0;
		9'd270: data = 5'd0;
		9'd271: data = 5'd0;
		9'd272: data = 5'd0;
		9'd273: data = 5'd0;
		9'd274: data = 5'd0;
		9'd275: data = 5'd0;
		9'd276: data = 5'd0;
		9'd277: data = 5'd0;
		9'd278: data = 5'd0;
		9'd279: data = 5'd3;
		9'd280: data = 5'd2;
		9'd281: data = 5'd4;
		9'd282: data = 5'd2;
		9'd283: data = 5'd0;
		9'd284: data = 5'd0;
		9'd285: data = 5'd0;
		9'd286: data = 5'd1;
		9'd287: data = 5'd7;
		9'd288: data = 5'd4;
		9'd289: data = 5'd0;
		9'd290: data = 5'd0;
		9'd291: data = 5'd0;
		9'd292: data = 5'd0;
		9'd293: data = 5'd0;
		9'd294: data = 5'd2;
		9'd295: data = 5'd0;
		9'd296: data = 5'd2;
		9'd297: data = 5'd0;
		9'd298: data = 5'd1;
		9'd299: data = 5'd0;
		9'd300: data = 5'd3;
		9'd301: data = 5'd0;
		9'd302: data = 5'd0;
		9'd303: data = 5'd1;
		9'd304: data = 5'd0;
		9'd305: data = 5'd0;
		9'd306: data = 5'd0;
		9'd307: data = 5'd0;
		9'd308: data = 5'd0;
		9'd309: data = 5'd5;
		9'd310: data = 5'd0;
		9'd311: data = 5'd0;
		9'd312: data = 5'd4;
		9'd313: data = 5'd6;
		9'd314: data = 5'd4;
		9'd315: data = 5'd0;
		9'd316: data = 5'd5;
		9'd317: data = 5'd3;
		9'd318: data = 5'd0;
		9'd319: data = 5'd0;
		9'd320: data = 5'd4;
		9'd321: data = 5'd0;
		9'd322: data = 5'd0;
		9'd323: data = 5'd0;
		9'd324: data = 5'd0;
		9'd325: data = 5'd0;
		9'd326: data = 5'd2;
		9'd327: data = 5'd5;
		9'd328: data = 5'd0;
		9'd329: data = 5'd0;
		9'd330: data = 5'd1;
		9'd331: data = 5'd0;
		9'd332: data = 5'd3;
		9'd333: data = 5'd0;
		9'd334: data = 5'd0;
		9'd335: data = 5'd3;
		9'd336: data = 5'd0;
		9'd337: data = 5'd0;
		9'd338: data = 5'd0;
		9'd339: data = 5'd0;
		9'd340: data = 5'd0;
		9'd341: data = 5'd5;
		9'd342: data = 5'd2;
		9'd343: data = 5'd4;
		9'd344: data = 5'd6;
		9'd345: data = 5'd0;
		9'd346: data = 5'd9;
		9'd347: data = 5'd0;
		9'd348: data = 5'd3;
		9'd349: data = 5'd0;
		9'd350: data = 5'd5;
		9'd351: data = 5'd2;
		9'd352: data = 5'd4;
		9'd353: data = 5'd16;
		9'd354: data = 5'd1;
		9'd355: data = 5'd0;
		9'd356: data = 5'd0;
		9'd357: data = 5'd0;
		9'd358: data = 5'd2;
		9'd359: data = 5'd3;
		9'd360: data = 5'd0;
		9'd361: data = 5'd0;
		9'd362: data = 5'd1;
		9'd363: data = 5'd0;
		9'd364: data = 5'd3;
		9'd365: data = 5'd0;
		9'd366: data = 5'd0;
		9'd367: data = 5'd0;
		9'd368: data = 5'd0;
		9'd369: data = 5'd0;
		9'd370: data = 5'd0;
		9'd371: data = 5'd0;
		9'd372: data = 5'd2;
		9'd373: data = 5'd1;
		9'd374: data = 5'd4;
		9'd375: data = 5'd6;
		9'd376: data = 5'd5;
		9'd377: data = 5'd0;
		9'd378: data = 5'd3;
		9'd379: data = 5'd5;
		9'd380: data = 5'd1;
		9'd381: data = 5'd2;
		9'd382: data = 5'd3;
		9'd383: data = 5'd4;
		9'd384: data = 5'd4;
		9'd385: data = 5'd17;
		9'd386: data = 5'd1;
		9'd387: data = 5'd0;
		9'd388: data = 5'd0;
		9'd389: data = 5'd0;
		9'd390: data = 5'd2;
		9'd391: data = 5'd3;
		9'd392: data = 5'd0;
		9'd393: data = 5'd0;
		9'd394: data = 5'd1;
		9'd395: data = 5'd0;
		9'd396: data = 5'd0;
		9'd397: data = 5'd0;
		9'd398: data = 5'd0;
		9'd399: data = 5'd0;
		9'd400: data = 5'd0;
		9'd401: data = 5'd0;
		9'd402: data = 5'd0;
		9'd403: data = 5'd5;
		9'd404: data = 5'd4;
		9'd405: data = 5'd4;
		9'd406: data = 5'd6;
		9'd407: data = 5'd0;
		9'd408: data = 5'd3;
		9'd409: data = 5'd0;
		9'd410: data = 5'd1;
		9'd411: data = 5'd0;
		9'd412: data = 5'd0;
		9'd413: data = 5'd4;
		9'd414: data = 5'd1;
		9'd415: data = 5'd6;
		9'd416: data = 5'd2;
		9'd417: data = 5'd18;
		9'd418: data = 5'd1;
		9'd419: data = 5'd0;
		9'd420: data = 5'd0;
		9'd421: data = 5'd0;
		9'd422: data = 5'd2;
		9'd423: data = 5'd3;
		9'd424: data = 5'd0;
		9'd425: data = 5'd0;
		9'd426: data = 5'd1;
		9'd427: data = 5'd0;
		9'd428: data = 5'd0;
		9'd429: data = 5'd6;
		9'd430: data = 5'd0;
		9'd431: data = 5'd0;
		9'd432: data = 5'd0;
		9'd433: data = 5'd0;
		9'd434: data = 5'd0;
		9'd435: data = 5'd1;
		9'd436: data = 5'd0;
		9'd437: data = 5'd0;
		9'd438: data = 5'd5;
		9'd439: data = 5'd0;
		9'd440: data = 5'd1;
		9'd441: data = 5'd5;
		9'd442: data = 5'd0;
		9'd443: data = 5'd4;
		9'd444: data = 5'd2;
		9'd445: data = 5'd6;
		9'd446: data = 5'd0;
		9'd447: data = 5'd0;
		9'd448: data = 5'd2;
		9'd449: data = 5'd19;
		9'd450: data = 5'd1;
		9'd451: data = 5'd0;
		9'd452: data = 5'd0;
		9'd453: data = 5'd0;
		9'd454: data = 5'd2;
		9'd455: data = 5'd3;
		9'd456: data = 5'd0;
		9'd457: data = 5'd0;
		9'd458: data = 5'd1;
		9'd459: data = 5'd0;
		9'd460: data = 5'd0;
		9'd461: data = 5'd2;
		9'd462: data = 5'd0;
		9'd463: data = 5'd0;
		9'd464: data = 5'd0;
		9'd465: data = 5'd0;
		9'd466: data = 5'd0;
		9'd467: data = 5'd6;
		9'd468: data = 5'd5;
		9'd469: data = 5'd0;
		9'd470: data = 5'd3;
		9'd471: data = 5'd0;
		9'd472: data = 5'd0;
		9'd473: data = 5'd1;
		9'd474: data = 5'd2;
		9'd475: data = 5'd6;
		9'd476: data = 5'd4;
		9'd477: data = 5'd0;
		9'd478: data = 5'd5;
		9'd479: data = 5'd5;
		9'd480: data = 5'd2;
		9'd481: data = 5'd11;
		9'd482: data = 5'd1;
		9'd483: data = 5'd0;
		9'd484: data = 5'd0;
		9'd485: data = 5'd0;
		9'd486: data = 5'd2;
		9'd487: data = 5'd5;
		9'd488: data = 5'd0;
		9'd489: data = 5'd0;
		9'd490: data = 5'd1;
		9'd491: data = 5'd0;
		9'd492: data = 5'd0;
		9'd493: data = 5'd0;
		9'd494: data = 5'd0;
		9'd495: data = 5'd0;
		9'd496: data = 5'd0;
		9'd497: data = 5'd5;
		9'd498: data = 5'd6;
		9'd499: data = 5'd0;
		9'd500: data = 5'd3;
		9'd501: data = 5'd0;
		9'd502: data = 5'd1;
		9'd503: data = 5'd0;
		9'd504: data = 5'd2;
		9'd505: data = 5'd2;
		9'd506: data = 5'd4;
		9'd507: data = 5'd6;
		9'd508: data = 5'd9;
		9'd509: data = 5'd0;
		9'd510: data = 5'd3;
		9'd511: data = 5'd1;
		default: data = 5'd0;
	endcase
end
endmodule

module layer1_N3_rsh_1(address, data);
input wire [8:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		9'd0: data = 1'd0;
		9'd1: data = 1'd0;
		9'd2: data = 1'd1;
		9'd3: data = 1'd1;
		9'd4: data = 1'd0;
		9'd5: data = 1'd1;
		9'd6: data = 1'd1;
		9'd7: data = 1'd1;
		9'd8: data = 1'd0;
		9'd9: data = 1'd1;
		9'd10: data = 1'd1;
		9'd11: data = 1'd1;
		9'd12: data = 1'd0;
		9'd13: data = 1'd1;
		9'd14: data = 1'd0;
		9'd15: data = 1'd1;
		9'd16: data = 1'd0;
		9'd17: data = 1'd0;
		9'd18: data = 1'd1;
		9'd19: data = 1'd1;
		9'd20: data = 1'd1;
		9'd21: data = 1'd1;
		9'd22: data = 1'd0;
		9'd23: data = 1'd1;
		9'd24: data = 1'd0;
		9'd25: data = 1'd1;
		9'd26: data = 1'd0;
		9'd27: data = 1'd0;
		9'd28: data = 1'd0;
		9'd29: data = 1'd0;
		9'd30: data = 1'd0;
		9'd31: data = 1'd0;
		9'd32: data = 1'd0;
		9'd33: data = 1'd0;
		9'd34: data = 1'd1;
		9'd35: data = 1'd1;
		9'd36: data = 1'd0;
		9'd37: data = 1'd1;
		9'd38: data = 1'd1;
		9'd39: data = 1'd1;
		9'd40: data = 1'd0;
		9'd41: data = 1'd1;
		9'd42: data = 1'd0;
		9'd43: data = 1'd1;
		9'd44: data = 1'd0;
		9'd45: data = 1'd1;
		9'd46: data = 1'd0;
		9'd47: data = 1'd1;
		9'd48: data = 1'd0;
		9'd49: data = 1'd0;
		9'd50: data = 1'd1;
		9'd51: data = 1'd1;
		9'd52: data = 1'd1;
		9'd53: data = 1'd1;
		9'd54: data = 1'd1;
		9'd55: data = 1'd1;
		9'd56: data = 1'd0;
		9'd57: data = 1'd1;
		9'd58: data = 1'd1;
		9'd59: data = 1'd0;
		9'd60: data = 1'd0;
		9'd61: data = 1'd0;
		9'd62: data = 1'd0;
		9'd63: data = 1'd0;
		9'd64: data = 1'd1;
		9'd65: data = 1'd0;
		9'd66: data = 1'd0;
		9'd67: data = 1'd1;
		9'd68: data = 1'd1;
		9'd69: data = 1'd1;
		9'd70: data = 1'd1;
		9'd71: data = 1'd1;
		9'd72: data = 1'd0;
		9'd73: data = 1'd1;
		9'd74: data = 1'd0;
		9'd75: data = 1'd1;
		9'd76: data = 1'd0;
		9'd77: data = 1'd1;
		9'd78: data = 1'd1;
		9'd79: data = 1'd1;
		9'd80: data = 1'd1;
		9'd81: data = 1'd1;
		9'd82: data = 1'd1;
		9'd83: data = 1'd1;
		9'd84: data = 1'd1;
		9'd85: data = 1'd1;
		9'd86: data = 1'd1;
		9'd87: data = 1'd1;
		9'd88: data = 1'd0;
		9'd89: data = 1'd1;
		9'd90: data = 1'd0;
		9'd91: data = 1'd1;
		9'd92: data = 1'd0;
		9'd93: data = 1'd0;
		9'd94: data = 1'd0;
		9'd95: data = 1'd0;
		9'd96: data = 1'd1;
		9'd97: data = 1'd1;
		9'd98: data = 1'd0;
		9'd99: data = 1'd1;
		9'd100: data = 1'd1;
		9'd101: data = 1'd1;
		9'd102: data = 1'd1;
		9'd103: data = 1'd1;
		9'd104: data = 1'd1;
		9'd105: data = 1'd1;
		9'd106: data = 1'd0;
		9'd107: data = 1'd1;
		9'd108: data = 1'd0;
		9'd109: data = 1'd1;
		9'd110: data = 1'd1;
		9'd111: data = 1'd1;
		9'd112: data = 1'd1;
		9'd113: data = 1'd1;
		9'd114: data = 1'd1;
		9'd115: data = 1'd1;
		9'd116: data = 1'd1;
		9'd117: data = 1'd1;
		9'd118: data = 1'd1;
		9'd119: data = 1'd1;
		9'd120: data = 1'd0;
		9'd121: data = 1'd1;
		9'd122: data = 1'd0;
		9'd123: data = 1'd1;
		9'd124: data = 1'd0;
		9'd125: data = 1'd0;
		9'd126: data = 1'd0;
		9'd127: data = 1'd0;
		9'd128: data = 1'd0;
		9'd129: data = 1'd1;
		9'd130: data = 1'd0;
		9'd131: data = 1'd1;
		9'd132: data = 1'd0;
		9'd133: data = 1'd1;
		9'd134: data = 1'd0;
		9'd135: data = 1'd1;
		9'd136: data = 1'd1;
		9'd137: data = 1'd1;
		9'd138: data = 1'd0;
		9'd139: data = 1'd1;
		9'd140: data = 1'd0;
		9'd141: data = 1'd1;
		9'd142: data = 1'd1;
		9'd143: data = 1'd1;
		9'd144: data = 1'd1;
		9'd145: data = 1'd1;
		9'd146: data = 1'd1;
		9'd147: data = 1'd1;
		9'd148: data = 1'd1;
		9'd149: data = 1'd1;
		9'd150: data = 1'd1;
		9'd151: data = 1'd1;
		9'd152: data = 1'd1;
		9'd153: data = 1'd1;
		9'd154: data = 1'd0;
		9'd155: data = 1'd1;
		9'd156: data = 1'd0;
		9'd157: data = 1'd0;
		9'd158: data = 1'd0;
		9'd159: data = 1'd0;
		9'd160: data = 1'd0;
		9'd161: data = 1'd1;
		9'd162: data = 1'd0;
		9'd163: data = 1'd1;
		9'd164: data = 1'd0;
		9'd165: data = 1'd1;
		9'd166: data = 1'd0;
		9'd167: data = 1'd1;
		9'd168: data = 1'd0;
		9'd169: data = 1'd1;
		9'd170: data = 1'd0;
		9'd171: data = 1'd1;
		9'd172: data = 1'd1;
		9'd173: data = 1'd1;
		9'd174: data = 1'd1;
		9'd175: data = 1'd1;
		9'd176: data = 1'd1;
		9'd177: data = 1'd1;
		9'd178: data = 1'd1;
		9'd179: data = 1'd1;
		9'd180: data = 1'd1;
		9'd181: data = 1'd1;
		9'd182: data = 1'd1;
		9'd183: data = 1'd1;
		9'd184: data = 1'd1;
		9'd185: data = 1'd1;
		9'd186: data = 1'd0;
		9'd187: data = 1'd0;
		9'd188: data = 1'd0;
		9'd189: data = 1'd0;
		9'd190: data = 1'd0;
		9'd191: data = 1'd0;
		9'd192: data = 1'd1;
		9'd193: data = 1'd1;
		9'd194: data = 1'd0;
		9'd195: data = 1'd1;
		9'd196: data = 1'd0;
		9'd197: data = 1'd1;
		9'd198: data = 1'd0;
		9'd199: data = 1'd1;
		9'd200: data = 1'd0;
		9'd201: data = 1'd1;
		9'd202: data = 1'd0;
		9'd203: data = 1'd1;
		9'd204: data = 1'd1;
		9'd205: data = 1'd1;
		9'd206: data = 1'd1;
		9'd207: data = 1'd0;
		9'd208: data = 1'd1;
		9'd209: data = 1'd1;
		9'd210: data = 1'd1;
		9'd211: data = 1'd1;
		9'd212: data = 1'd1;
		9'd213: data = 1'd1;
		9'd214: data = 1'd1;
		9'd215: data = 1'd1;
		9'd216: data = 1'd1;
		9'd217: data = 1'd1;
		9'd218: data = 1'd0;
		9'd219: data = 1'd0;
		9'd220: data = 1'd0;
		9'd221: data = 1'd0;
		9'd222: data = 1'd0;
		9'd223: data = 1'd0;
		9'd224: data = 1'd1;
		9'd225: data = 1'd1;
		9'd226: data = 1'd0;
		9'd227: data = 1'd1;
		9'd228: data = 1'd0;
		9'd229: data = 1'd1;
		9'd230: data = 1'd0;
		9'd231: data = 1'd1;
		9'd232: data = 1'd0;
		9'd233: data = 1'd1;
		9'd234: data = 1'd0;
		9'd235: data = 1'd1;
		9'd236: data = 1'd1;
		9'd237: data = 1'd1;
		9'd238: data = 1'd1;
		9'd239: data = 1'd0;
		9'd240: data = 1'd1;
		9'd241: data = 1'd1;
		9'd242: data = 1'd1;
		9'd243: data = 1'd1;
		9'd244: data = 1'd1;
		9'd245: data = 1'd1;
		9'd246: data = 1'd0;
		9'd247: data = 1'd1;
		9'd248: data = 1'd0;
		9'd249: data = 1'd0;
		9'd250: data = 1'd0;
		9'd251: data = 1'd0;
		9'd252: data = 1'd0;
		9'd253: data = 1'd0;
		9'd254: data = 1'd0;
		9'd255: data = 1'd0;
		9'd256: data = 1'd0;
		9'd257: data = 1'd1;
		9'd258: data = 1'd0;
		9'd259: data = 1'd1;
		9'd260: data = 1'd0;
		9'd261: data = 1'd1;
		9'd262: data = 1'd0;
		9'd263: data = 1'd1;
		9'd264: data = 1'd0;
		9'd265: data = 1'd1;
		9'd266: data = 1'd0;
		9'd267: data = 1'd1;
		9'd268: data = 1'd1;
		9'd269: data = 1'd1;
		9'd270: data = 1'd1;
		9'd271: data = 1'd0;
		9'd272: data = 1'd1;
		9'd273: data = 1'd1;
		9'd274: data = 1'd1;
		9'd275: data = 1'd1;
		9'd276: data = 1'd0;
		9'd277: data = 1'd1;
		9'd278: data = 1'd0;
		9'd279: data = 1'd1;
		9'd280: data = 1'd0;
		9'd281: data = 1'd0;
		9'd282: data = 1'd0;
		9'd283: data = 1'd1;
		9'd284: data = 1'd0;
		9'd285: data = 1'd1;
		9'd286: data = 1'd0;
		9'd287: data = 1'd0;
		9'd288: data = 1'd0;
		9'd289: data = 1'd1;
		9'd290: data = 1'd0;
		9'd291: data = 1'd1;
		9'd292: data = 1'd0;
		9'd293: data = 1'd1;
		9'd294: data = 1'd0;
		9'd295: data = 1'd1;
		9'd296: data = 1'd0;
		9'd297: data = 1'd1;
		9'd298: data = 1'd1;
		9'd299: data = 1'd1;
		9'd300: data = 1'd1;
		9'd301: data = 1'd1;
		9'd302: data = 1'd1;
		9'd303: data = 1'd1;
		9'd304: data = 1'd1;
		9'd305: data = 1'd1;
		9'd306: data = 1'd1;
		9'd307: data = 1'd1;
		9'd308: data = 1'd0;
		9'd309: data = 1'd1;
		9'd310: data = 1'd0;
		9'd311: data = 1'd0;
		9'd312: data = 1'd0;
		9'd313: data = 1'd0;
		9'd314: data = 1'd0;
		9'd315: data = 1'd1;
		9'd316: data = 1'd0;
		9'd317: data = 1'd1;
		9'd318: data = 1'd0;
		9'd319: data = 1'd0;
		9'd320: data = 1'd0;
		9'd321: data = 1'd1;
		9'd322: data = 1'd0;
		9'd323: data = 1'd1;
		9'd324: data = 1'd0;
		9'd325: data = 1'd1;
		9'd326: data = 1'd0;
		9'd327: data = 1'd1;
		9'd328: data = 1'd0;
		9'd329: data = 1'd1;
		9'd330: data = 1'd1;
		9'd331: data = 1'd1;
		9'd332: data = 1'd1;
		9'd333: data = 1'd1;
		9'd334: data = 1'd1;
		9'd335: data = 1'd1;
		9'd336: data = 1'd1;
		9'd337: data = 1'd1;
		9'd338: data = 1'd1;
		9'd339: data = 1'd1;
		9'd340: data = 1'd0;
		9'd341: data = 1'd1;
		9'd342: data = 1'd0;
		9'd343: data = 1'd0;
		9'd344: data = 1'd0;
		9'd345: data = 1'd1;
		9'd346: data = 1'd0;
		9'd347: data = 1'd1;
		9'd348: data = 1'd0;
		9'd349: data = 1'd0;
		9'd350: data = 1'd0;
		9'd351: data = 1'd0;
		9'd352: data = 1'd0;
		9'd353: data = 1'd0;
		9'd354: data = 1'd1;
		9'd355: data = 1'd1;
		9'd356: data = 1'd0;
		9'd357: data = 1'd1;
		9'd358: data = 1'd0;
		9'd359: data = 1'd1;
		9'd360: data = 1'd0;
		9'd361: data = 1'd1;
		9'd362: data = 1'd1;
		9'd363: data = 1'd1;
		9'd364: data = 1'd1;
		9'd365: data = 1'd1;
		9'd366: data = 1'd1;
		9'd367: data = 1'd1;
		9'd368: data = 1'd1;
		9'd369: data = 1'd1;
		9'd370: data = 1'd1;
		9'd371: data = 1'd1;
		9'd372: data = 1'd0;
		9'd373: data = 1'd1;
		9'd374: data = 1'd0;
		9'd375: data = 1'd0;
		9'd376: data = 1'd1;
		9'd377: data = 1'd1;
		9'd378: data = 1'd1;
		9'd379: data = 1'd1;
		9'd380: data = 1'd0;
		9'd381: data = 1'd0;
		9'd382: data = 1'd0;
		9'd383: data = 1'd0;
		9'd384: data = 1'd0;
		9'd385: data = 1'd0;
		9'd386: data = 1'd1;
		9'd387: data = 1'd1;
		9'd388: data = 1'd0;
		9'd389: data = 1'd1;
		9'd390: data = 1'd0;
		9'd391: data = 1'd1;
		9'd392: data = 1'd0;
		9'd393: data = 1'd1;
		9'd394: data = 1'd1;
		9'd395: data = 1'd1;
		9'd396: data = 1'd1;
		9'd397: data = 1'd1;
		9'd398: data = 1'd1;
		9'd399: data = 1'd1;
		9'd400: data = 1'd1;
		9'd401: data = 1'd1;
		9'd402: data = 1'd1;
		9'd403: data = 1'd1;
		9'd404: data = 1'd0;
		9'd405: data = 1'd0;
		9'd406: data = 1'd0;
		9'd407: data = 1'd1;
		9'd408: data = 1'd1;
		9'd409: data = 1'd1;
		9'd410: data = 1'd1;
		9'd411: data = 1'd0;
		9'd412: data = 1'd0;
		9'd413: data = 1'd0;
		9'd414: data = 1'd0;
		9'd415: data = 1'd0;
		9'd416: data = 1'd0;
		9'd417: data = 1'd0;
		9'd418: data = 1'd1;
		9'd419: data = 1'd1;
		9'd420: data = 1'd0;
		9'd421: data = 1'd1;
		9'd422: data = 1'd0;
		9'd423: data = 1'd1;
		9'd424: data = 1'd0;
		9'd425: data = 1'd1;
		9'd426: data = 1'd1;
		9'd427: data = 1'd1;
		9'd428: data = 1'd1;
		9'd429: data = 1'd0;
		9'd430: data = 1'd1;
		9'd431: data = 1'd1;
		9'd432: data = 1'd1;
		9'd433: data = 1'd1;
		9'd434: data = 1'd1;
		9'd435: data = 1'd1;
		9'd436: data = 1'd1;
		9'd437: data = 1'd1;
		9'd438: data = 1'd1;
		9'd439: data = 1'd1;
		9'd440: data = 1'd1;
		9'd441: data = 1'd1;
		9'd442: data = 1'd0;
		9'd443: data = 1'd0;
		9'd444: data = 1'd0;
		9'd445: data = 1'd0;
		9'd446: data = 1'd0;
		9'd447: data = 1'd1;
		9'd448: data = 1'd0;
		9'd449: data = 1'd0;
		9'd450: data = 1'd1;
		9'd451: data = 1'd1;
		9'd452: data = 1'd0;
		9'd453: data = 1'd1;
		9'd454: data = 1'd0;
		9'd455: data = 1'd1;
		9'd456: data = 1'd0;
		9'd457: data = 1'd1;
		9'd458: data = 1'd1;
		9'd459: data = 1'd1;
		9'd460: data = 1'd1;
		9'd461: data = 1'd0;
		9'd462: data = 1'd1;
		9'd463: data = 1'd1;
		9'd464: data = 1'd1;
		9'd465: data = 1'd1;
		9'd466: data = 1'd1;
		9'd467: data = 1'd0;
		9'd468: data = 1'd1;
		9'd469: data = 1'd1;
		9'd470: data = 1'd1;
		9'd471: data = 1'd1;
		9'd472: data = 1'd0;
		9'd473: data = 1'd1;
		9'd474: data = 1'd0;
		9'd475: data = 1'd0;
		9'd476: data = 1'd0;
		9'd477: data = 1'd1;
		9'd478: data = 1'd0;
		9'd479: data = 1'd1;
		9'd480: data = 1'd0;
		9'd481: data = 1'd0;
		9'd482: data = 1'd1;
		9'd483: data = 1'd1;
		9'd484: data = 1'd0;
		9'd485: data = 1'd1;
		9'd486: data = 1'd0;
		9'd487: data = 1'd1;
		9'd488: data = 1'd0;
		9'd489: data = 1'd1;
		9'd490: data = 1'd1;
		9'd491: data = 1'd1;
		9'd492: data = 1'd1;
		9'd493: data = 1'd0;
		9'd494: data = 1'd1;
		9'd495: data = 1'd1;
		9'd496: data = 1'd1;
		9'd497: data = 1'd1;
		9'd498: data = 1'd0;
		9'd499: data = 1'd1;
		9'd500: data = 1'd1;
		9'd501: data = 1'd1;
		9'd502: data = 1'd1;
		9'd503: data = 1'd1;
		9'd504: data = 1'd0;
		9'd505: data = 1'd0;
		9'd506: data = 1'd0;
		9'd507: data = 1'd0;
		9'd508: data = 1'd0;
		9'd509: data = 1'd1;
		9'd510: data = 1'd0;
		9'd511: data = 1'd1;
		default: data = 1'd0;
	endcase
end
endmodule

module layer1_N3(address, data);
input wire [11:0] address;
output reg [3:0] data;

wire [4:0] i; layer1_N3_idx_1 idx_1_inst(address[11:3], i);
wire [0:0] t; layer1_N3_rsh_1 rsh_1_inst(address[11:3], t);
wire [3:0] b; layer1_N3_2 layer1_N3_2_inst(address[11:3], b);
wire [1:0] u; layer1_N3_ust_1 ust_1_inst({i, address[2:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule
