module layer0 (input [63:0] address, output [127:0] data);

wire [11:0] layer0_N0_wire = {address[15], address[14], address[13], address[12], address[35], address[34], address[33], address[32], address[55], address[54], address[53], address[52]};
layer0_N0 layer0_N0_inst (.address(layer0_N0_wire), .data(data[3:0]));

wire [11:0] layer0_N1_wire = {address[19], address[18], address[17], address[16], address[43], address[42], address[41], address[40], address[63], address[62], address[61], address[60]};
layer0_N1 layer0_N1_inst (.address(layer0_N1_wire), .data(data[7:4]));

wire [11:0] layer0_N2_wire = {address[7], address[6], address[5], address[4], address[39], address[38], address[37], address[36], address[59], address[58], address[57], address[56]};
layer0_N2 layer0_N2_inst (.address(layer0_N2_wire), .data(data[11:8]));

wire [11:0] layer0_N3_wire = {address[27], address[26], address[25], address[24], address[39], address[38], address[37], address[36], address[51], address[50], address[49], address[48]};
layer0_N3 layer0_N3_inst (.address(layer0_N3_wire), .data(data[15:12]));

wire [11:0] layer0_N4_wire = {address[7], address[6], address[5], address[4], address[51], address[50], address[49], address[48], address[63], address[62], address[61], address[60]};
layer0_N4 layer0_N4_inst (.address(layer0_N4_wire), .data(data[19:16]));

wire [11:0] layer0_N5_wire = {address[47], address[46], address[45], address[44], address[51], address[50], address[49], address[48], address[63], address[62], address[61], address[60]};
layer0_N5 layer0_N5_inst (.address(layer0_N5_wire), .data(data[23:20]));

wire [11:0] layer0_N6_wire = {address[15], address[14], address[13], address[12], address[35], address[34], address[33], address[32], address[51], address[50], address[49], address[48]};
layer0_N6 layer0_N6_inst (.address(layer0_N6_wire), .data(data[27:24]));

wire [11:0] layer0_N7_wire = {address[15], address[14], address[13], address[12], address[19], address[18], address[17], address[16], address[51], address[50], address[49], address[48]};
layer0_N7 layer0_N7_inst (.address(layer0_N7_wire), .data(data[31:28]));

wire [11:0] layer0_N8_wire = {address[43], address[42], address[41], address[40], address[51], address[50], address[49], address[48], address[59], address[58], address[57], address[56]};
layer0_N8 layer0_N8_inst (.address(layer0_N8_wire), .data(data[35:32]));

wire [11:0] layer0_N9_wire = {address[23], address[22], address[21], address[20], address[35], address[34], address[33], address[32], address[51], address[50], address[49], address[48]};
layer0_N9 layer0_N9_inst (.address(layer0_N9_wire), .data(data[39:36]));

wire [11:0] layer0_N10_wire = {address[23], address[22], address[21], address[20], address[39], address[38], address[37], address[36], address[43], address[42], address[41], address[40]};
layer0_N10 layer0_N10_inst (.address(layer0_N10_wire), .data(data[43:40]));

wire [11:0] layer0_N11_wire = {address[11], address[10], address[9], address[8], address[23], address[22], address[21], address[20], address[59], address[58], address[57], address[56]};
layer0_N11 layer0_N11_inst (.address(layer0_N11_wire), .data(data[47:44]));

wire [11:0] layer0_N12_wire = {address[3], address[2], address[1], address[0], address[19], address[18], address[17], address[16], address[27], address[26], address[25], address[24]};
layer0_N12 layer0_N12_inst (.address(layer0_N12_wire), .data(data[51:48]));

wire [11:0] layer0_N13_wire = {address[27], address[26], address[25], address[24], address[39], address[38], address[37], address[36], address[55], address[54], address[53], address[52]};
layer0_N13 layer0_N13_inst (.address(layer0_N13_wire), .data(data[55:52]));

wire [11:0] layer0_N14_wire = {address[7], address[6], address[5], address[4], address[19], address[18], address[17], address[16], address[51], address[50], address[49], address[48]};
layer0_N14 layer0_N14_inst (.address(layer0_N14_wire), .data(data[59:56]));

wire [11:0] layer0_N15_wire = {address[31], address[30], address[29], address[28], address[47], address[46], address[45], address[44], address[55], address[54], address[53], address[52]};
layer0_N15 layer0_N15_inst (.address(layer0_N15_wire), .data(data[63:60]));

wire [11:0] layer0_N16_wire = {address[3], address[2], address[1], address[0], address[15], address[14], address[13], address[12], address[31], address[30], address[29], address[28]};
layer0_N16 layer0_N16_inst (.address(layer0_N16_wire), .data(data[67:64]));

wire [11:0] layer0_N17_wire = {address[47], address[46], address[45], address[44], address[55], address[54], address[53], address[52], address[59], address[58], address[57], address[56]};
layer0_N17 layer0_N17_inst (.address(layer0_N17_wire), .data(data[71:68]));

wire [11:0] layer0_N18_wire = {address[11], address[10], address[9], address[8], address[27], address[26], address[25], address[24], address[43], address[42], address[41], address[40]};
layer0_N18 layer0_N18_inst (.address(layer0_N18_wire), .data(data[75:72]));

wire [11:0] layer0_N19_wire = {address[23], address[22], address[21], address[20], address[43], address[42], address[41], address[40], address[51], address[50], address[49], address[48]};
layer0_N19 layer0_N19_inst (.address(layer0_N19_wire), .data(data[79:76]));

wire [11:0] layer0_N20_wire = {address[3], address[2], address[1], address[0], address[19], address[18], address[17], address[16], address[51], address[50], address[49], address[48]};
layer0_N20 layer0_N20_inst (.address(layer0_N20_wire), .data(data[83:80]));

wire [11:0] layer0_N21_wire = {address[35], address[34], address[33], address[32], address[55], address[54], address[53], address[52], address[59], address[58], address[57], address[56]};
layer0_N21 layer0_N21_inst (.address(layer0_N21_wire), .data(data[87:84]));

wire [11:0] layer0_N22_wire = {address[27], address[26], address[25], address[24], address[35], address[34], address[33], address[32], address[39], address[38], address[37], address[36]};
layer0_N22 layer0_N22_inst (.address(layer0_N22_wire), .data(data[91:88]));

wire [11:0] layer0_N23_wire = {address[3], address[2], address[1], address[0], address[11], address[10], address[9], address[8], address[55], address[54], address[53], address[52]};
layer0_N23 layer0_N23_inst (.address(layer0_N23_wire), .data(data[95:92]));

wire [11:0] layer0_N24_wire = {address[15], address[14], address[13], address[12], address[19], address[18], address[17], address[16], address[27], address[26], address[25], address[24]};
layer0_N24 layer0_N24_inst (.address(layer0_N24_wire), .data(data[99:96]));

wire [11:0] layer0_N25_wire = {address[15], address[14], address[13], address[12], address[31], address[30], address[29], address[28], address[59], address[58], address[57], address[56]};
layer0_N25 layer0_N25_inst (.address(layer0_N25_wire), .data(data[103:100]));

wire [11:0] layer0_N26_wire = {address[31], address[30], address[29], address[28], address[35], address[34], address[33], address[32], address[63], address[62], address[61], address[60]};
layer0_N26 layer0_N26_inst (.address(layer0_N26_wire), .data(data[107:104]));

wire [11:0] layer0_N27_wire = {address[3], address[2], address[1], address[0], address[15], address[14], address[13], address[12], address[51], address[50], address[49], address[48]};
layer0_N27 layer0_N27_inst (.address(layer0_N27_wire), .data(data[111:108]));

wire [11:0] layer0_N28_wire = {address[7], address[6], address[5], address[4], address[19], address[18], address[17], address[16], address[31], address[30], address[29], address[28]};
layer0_N28 layer0_N28_inst (.address(layer0_N28_wire), .data(data[115:112]));

wire [11:0] layer0_N29_wire = {address[3], address[2], address[1], address[0], address[11], address[10], address[9], address[8], address[27], address[26], address[25], address[24]};
layer0_N29 layer0_N29_inst (.address(layer0_N29_wire), .data(data[119:116]));

wire [11:0] layer0_N30_wire = {address[3], address[2], address[1], address[0], address[19], address[18], address[17], address[16], address[47], address[46], address[45], address[44]};
layer0_N30 layer0_N30_inst (.address(layer0_N30_wire), .data(data[123:120]));

wire [11:0] layer0_N31_wire = {address[11], address[10], address[9], address[8], address[23], address[22], address[21], address[20], address[31], address[30], address[29], address[28]};
layer0_N31 layer0_N31_inst (.address(layer0_N31_wire), .data(data[127:124]));

endmodule