
module layer1_N4_ust_3(address, data);
input wire [3:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		4'd0: data = 1'd1;
		4'd1: data = 1'd0;
		4'd2: data = 1'd0;
		4'd3: data = 1'd0;
		4'd4: data = 1'd1;
		4'd5: data = 1'd0;
		4'd6: data = 1'd0;
		4'd7: data = 1'd0;
		4'd8: data = 1'd1;
		4'd9: data = 1'd1;
		4'd10: data = 1'd0;
		4'd11: data = 1'd0;
		4'd12: data = 1'd1;
		4'd13: data = 1'd1;
		4'd14: data = 1'd0;
		4'd15: data = 1'd0;
		default: data = 1'd0;
	endcase
end
endmodule

module layer1_N4_idx_3(address, data);
input wire [2:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		3'd0: data = 1'd0;
		3'd1: data = 1'd0;
		3'd2: data = 1'd0;
		3'd3: data = 1'd0;
		3'd4: data = 1'd0;
		3'd5: data = 1'd0;
		3'd6: data = 1'd0;
		3'd7: data = 1'd1;
		default: data = 1'd0;
	endcase
end
endmodule

module layer1_N4_rsh_3(address, data);
input wire [2:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		3'd0: data = 1'd1;
		3'd1: data = 1'd1;
		3'd2: data = 1'd1;
		3'd3: data = 1'd1;
		3'd4: data = 1'd0;
		3'd5: data = 1'd0;
		3'd6: data = 1'd0;
		3'd7: data = 1'd0;
		default: data = 1'd0;
	endcase
end
endmodule

module layer1_N4_3(address, data);
input wire [5:0] address;
output reg [0:0] data;

wire [0:0] i; layer1_N4_idx_3 idx_3_inst(address[5:3], i);
wire [0:0] t; layer1_N4_rsh_3 rsh_3_inst(address[5:3], t);
wire [0:0] u; layer1_N4_ust_3 ust_3_inst({i, address[2:0]}, u);

always @(*) begin
	data = (u >> t);
end
endmodule

module layer1_N4_ust_2(address, data);
input wire [8:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		9'd0: data = 1'd1;
		9'd1: data = 1'd1;
		9'd2: data = 1'd1;
		9'd3: data = 1'd0;
		9'd4: data = 1'd1;
		9'd5: data = 1'd1;
		9'd6: data = 1'd1;
		9'd7: data = 1'd0;
		9'd8: data = 1'd1;
		9'd9: data = 1'd1;
		9'd10: data = 1'd1;
		9'd11: data = 1'd0;
		9'd12: data = 1'd1;
		9'd13: data = 1'd1;
		9'd14: data = 1'd1;
		9'd15: data = 1'd0;
		9'd16: data = 1'd0;
		9'd17: data = 1'd0;
		9'd18: data = 1'd1;
		9'd19: data = 1'd0;
		9'd20: data = 1'd0;
		9'd21: data = 1'd0;
		9'd22: data = 1'd1;
		9'd23: data = 1'd0;
		9'd24: data = 1'd0;
		9'd25: data = 1'd0;
		9'd26: data = 1'd1;
		9'd27: data = 1'd0;
		9'd28: data = 1'd0;
		9'd29: data = 1'd0;
		9'd30: data = 1'd1;
		9'd31: data = 1'd0;
		9'd32: data = 1'd1;
		9'd33: data = 1'd1;
		9'd34: data = 1'd1;
		9'd35: data = 1'd1;
		9'd36: data = 1'd1;
		9'd37: data = 1'd1;
		9'd38: data = 1'd1;
		9'd39: data = 1'd1;
		9'd40: data = 1'd1;
		9'd41: data = 1'd1;
		9'd42: data = 1'd1;
		9'd43: data = 1'd1;
		9'd44: data = 1'd1;
		9'd45: data = 1'd1;
		9'd46: data = 1'd1;
		9'd47: data = 1'd0;
		9'd48: data = 1'd1;
		9'd49: data = 1'd1;
		9'd50: data = 1'd1;
		9'd51: data = 1'd1;
		9'd52: data = 1'd1;
		9'd53: data = 1'd1;
		9'd54: data = 1'd1;
		9'd55: data = 1'd0;
		9'd56: data = 1'd1;
		9'd57: data = 1'd1;
		9'd58: data = 1'd1;
		9'd59: data = 1'd0;
		9'd60: data = 1'd1;
		9'd61: data = 1'd1;
		9'd62: data = 1'd1;
		9'd63: data = 1'd0;
		9'd64: data = 1'd1;
		9'd65: data = 1'd1;
		9'd66: data = 1'd1;
		9'd67: data = 1'd1;
		9'd68: data = 1'd1;
		9'd69: data = 1'd1;
		9'd70: data = 1'd1;
		9'd71: data = 1'd1;
		9'd72: data = 1'd1;
		9'd73: data = 1'd1;
		9'd74: data = 1'd1;
		9'd75: data = 1'd0;
		9'd76: data = 1'd1;
		9'd77: data = 1'd1;
		9'd78: data = 1'd1;
		9'd79: data = 1'd0;
		9'd80: data = 1'd1;
		9'd81: data = 1'd1;
		9'd82: data = 1'd1;
		9'd83: data = 1'd0;
		9'd84: data = 1'd0;
		9'd85: data = 1'd0;
		9'd86: data = 1'd0;
		9'd87: data = 1'd0;
		9'd88: data = 1'd0;
		9'd89: data = 1'd0;
		9'd90: data = 1'd0;
		9'd91: data = 1'd0;
		9'd92: data = 1'd0;
		9'd93: data = 1'd0;
		9'd94: data = 1'd0;
		9'd95: data = 1'd0;
		9'd96: data = 1'd0;
		9'd97: data = 1'd1;
		9'd98: data = 1'd1;
		9'd99: data = 1'd0;
		9'd100: data = 1'd0;
		9'd101: data = 1'd1;
		9'd102: data = 1'd1;
		9'd103: data = 1'd0;
		9'd104: data = 1'd0;
		9'd105: data = 1'd0;
		9'd106: data = 1'd1;
		9'd107: data = 1'd0;
		9'd108: data = 1'd0;
		9'd109: data = 1'd0;
		9'd110: data = 1'd1;
		9'd111: data = 1'd0;
		9'd112: data = 1'd1;
		9'd113: data = 1'd1;
		9'd114: data = 1'd1;
		9'd115: data = 1'd0;
		9'd116: data = 1'd1;
		9'd117: data = 1'd1;
		9'd118: data = 1'd1;
		9'd119: data = 1'd0;
		9'd120: data = 1'd1;
		9'd121: data = 1'd1;
		9'd122: data = 1'd1;
		9'd123: data = 1'd0;
		9'd124: data = 1'd0;
		9'd125: data = 1'd1;
		9'd126: data = 1'd1;
		9'd127: data = 1'd0;
		9'd128: data = 1'd1;
		9'd129: data = 1'd1;
		9'd130: data = 1'd1;
		9'd131: data = 1'd0;
		9'd132: data = 1'd1;
		9'd133: data = 1'd1;
		9'd134: data = 1'd1;
		9'd135: data = 1'd0;
		9'd136: data = 1'd1;
		9'd137: data = 1'd1;
		9'd138: data = 1'd1;
		9'd139: data = 1'd0;
		9'd140: data = 1'd1;
		9'd141: data = 1'd1;
		9'd142: data = 1'd0;
		9'd143: data = 1'd0;
		9'd144: data = 1'd1;
		9'd145: data = 1'd0;
		9'd146: data = 1'd0;
		9'd147: data = 1'd0;
		9'd148: data = 1'd0;
		9'd149: data = 1'd0;
		9'd150: data = 1'd0;
		9'd151: data = 1'd0;
		9'd152: data = 1'd0;
		9'd153: data = 1'd0;
		9'd154: data = 1'd0;
		9'd155: data = 1'd0;
		9'd156: data = 1'd0;
		9'd157: data = 1'd0;
		9'd158: data = 1'd0;
		9'd159: data = 1'd0;
		9'd160: data = 1'd1;
		9'd161: data = 1'd1;
		9'd162: data = 1'd1;
		9'd163: data = 1'd0;
		9'd164: data = 1'd0;
		9'd165: data = 1'd0;
		9'd166: data = 1'd1;
		9'd167: data = 1'd0;
		9'd168: data = 1'd0;
		9'd169: data = 1'd0;
		9'd170: data = 1'd0;
		9'd171: data = 1'd0;
		9'd172: data = 1'd0;
		9'd173: data = 1'd0;
		9'd174: data = 1'd0;
		9'd175: data = 1'd0;
		9'd176: data = 1'd1;
		9'd177: data = 1'd1;
		9'd178: data = 1'd1;
		9'd179: data = 1'd0;
		9'd180: data = 1'd0;
		9'd181: data = 1'd1;
		9'd182: data = 1'd1;
		9'd183: data = 1'd0;
		9'd184: data = 1'd0;
		9'd185: data = 1'd0;
		9'd186: data = 1'd0;
		9'd187: data = 1'd0;
		9'd188: data = 1'd0;
		9'd189: data = 1'd0;
		9'd190: data = 1'd0;
		9'd191: data = 1'd0;
		9'd192: data = 1'd1;
		9'd193: data = 1'd1;
		9'd194: data = 1'd1;
		9'd195: data = 1'd0;
		9'd196: data = 1'd1;
		9'd197: data = 1'd1;
		9'd198: data = 1'd1;
		9'd199: data = 1'd0;
		9'd200: data = 1'd0;
		9'd201: data = 1'd1;
		9'd202: data = 1'd0;
		9'd203: data = 1'd0;
		9'd204: data = 1'd0;
		9'd205: data = 1'd0;
		9'd206: data = 1'd0;
		9'd207: data = 1'd0;
		9'd208: data = 1'd0;
		9'd209: data = 1'd0;
		9'd210: data = 1'd0;
		9'd211: data = 1'd0;
		9'd212: data = 1'd0;
		9'd213: data = 1'd0;
		9'd214: data = 1'd0;
		9'd215: data = 1'd0;
		9'd216: data = 1'd0;
		9'd217: data = 1'd0;
		9'd218: data = 1'd0;
		9'd219: data = 1'd0;
		9'd220: data = 1'd0;
		9'd221: data = 1'd0;
		9'd222: data = 1'd1;
		9'd223: data = 1'd0;
		9'd224: data = 1'd1;
		9'd225: data = 1'd1;
		9'd226: data = 1'd1;
		9'd227: data = 1'd0;
		9'd228: data = 1'd1;
		9'd229: data = 1'd1;
		9'd230: data = 1'd1;
		9'd231: data = 1'd0;
		9'd232: data = 1'd0;
		9'd233: data = 1'd1;
		9'd234: data = 1'd1;
		9'd235: data = 1'd0;
		9'd236: data = 1'd0;
		9'd237: data = 1'd0;
		9'd238: data = 1'd1;
		9'd239: data = 1'd0;
		9'd240: data = 1'd0;
		9'd241: data = 1'd0;
		9'd242: data = 1'd1;
		9'd243: data = 1'd0;
		9'd244: data = 1'd0;
		9'd245: data = 1'd0;
		9'd246: data = 1'd0;
		9'd247: data = 1'd0;
		9'd248: data = 1'd0;
		9'd249: data = 1'd0;
		9'd250: data = 1'd1;
		9'd251: data = 1'd0;
		9'd252: data = 1'd0;
		9'd253: data = 1'd0;
		9'd254: data = 1'd1;
		9'd255: data = 1'd0;
		9'd256: data = 1'd1;
		9'd257: data = 1'd1;
		9'd258: data = 1'd1;
		9'd259: data = 1'd0;
		9'd260: data = 1'd1;
		9'd261: data = 1'd1;
		9'd262: data = 1'd1;
		9'd263: data = 1'd0;
		9'd264: data = 1'd0;
		9'd265: data = 1'd1;
		9'd266: data = 1'd1;
		9'd267: data = 1'd0;
		9'd268: data = 1'd0;
		9'd269: data = 1'd1;
		9'd270: data = 1'd1;
		9'd271: data = 1'd0;
		9'd272: data = 1'd0;
		9'd273: data = 1'd1;
		9'd274: data = 1'd1;
		9'd275: data = 1'd0;
		9'd276: data = 1'd0;
		9'd277: data = 1'd1;
		9'd278: data = 1'd1;
		9'd279: data = 1'd0;
		9'd280: data = 1'd0;
		9'd281: data = 1'd1;
		9'd282: data = 1'd1;
		9'd283: data = 1'd0;
		9'd284: data = 1'd0;
		9'd285: data = 1'd0;
		9'd286: data = 1'd1;
		9'd287: data = 1'd0;
		9'd288: data = 1'd1;
		9'd289: data = 1'd1;
		9'd290: data = 1'd1;
		9'd291: data = 1'd0;
		9'd292: data = 1'd0;
		9'd293: data = 1'd1;
		9'd294: data = 1'd1;
		9'd295: data = 1'd0;
		9'd296: data = 1'd0;
		9'd297: data = 1'd1;
		9'd298: data = 1'd1;
		9'd299: data = 1'd0;
		9'd300: data = 1'd0;
		9'd301: data = 1'd1;
		9'd302: data = 1'd1;
		9'd303: data = 1'd0;
		default: data = 1'd0;
	endcase
end
endmodule

module layer1_N4_idx_2(address, data);
input wire [5:0] address;
output reg [4:0] data;

always @(*) begin
	case(address)
		6'd0: data = 5'd8;
		6'd1: data = 5'd0;
		6'd2: data = 5'd0;
		6'd3: data = 5'd0;
		6'd4: data = 5'd0;
		6'd5: data = 5'd0;
		6'd6: data = 5'd0;
		6'd7: data = 5'd0;
		6'd8: data = 5'd3;
		6'd9: data = 5'd9;
		6'd10: data = 5'd0;
		6'd11: data = 5'd0;
		6'd12: data = 5'd4;
		6'd13: data = 5'd5;
		6'd14: data = 5'd0;
		6'd15: data = 5'd0;
		6'd16: data = 5'd2;
		6'd17: data = 5'd5;
		6'd18: data = 5'd0;
		6'd19: data = 5'd0;
		6'd20: data = 5'd2;
		6'd21: data = 5'd10;
		6'd22: data = 5'd0;
		6'd23: data = 5'd0;
		6'd24: data = 5'd2;
		6'd25: data = 5'd11;
		6'd26: data = 5'd0;
		6'd27: data = 5'd0;
		6'd28: data = 5'd2;
		6'd29: data = 5'd12;
		6'd30: data = 5'd13;
		6'd31: data = 5'd1;
		6'd32: data = 5'd0;
		6'd33: data = 5'd14;
		6'd34: data = 5'd15;
		6'd35: data = 5'd1;
		6'd36: data = 5'd0;
		6'd37: data = 5'd16;
		6'd38: data = 5'd6;
		6'd39: data = 5'd1;
		6'd40: data = 5'd0;
		6'd41: data = 5'd7;
		6'd42: data = 5'd6;
		6'd43: data = 5'd1;
		6'd44: data = 5'd0;
		6'd45: data = 5'd7;
		6'd46: data = 5'd17;
		6'd47: data = 5'd1;
		6'd48: data = 5'd0;
		6'd49: data = 5'd0;
		6'd50: data = 5'd18;
		6'd51: data = 5'd1;
		6'd52: data = 5'd0;
		6'd53: data = 5'd4;
		6'd54: data = 5'd0;
		6'd55: data = 5'd0;
		6'd56: data = 5'd0;
		6'd57: data = 5'd0;
		6'd58: data = 5'd0;
		6'd59: data = 5'd0;
		6'd60: data = 5'd0;
		6'd61: data = 5'd0;
		6'd62: data = 5'd3;
		6'd63: data = 5'd0;
		default: data = 5'd0;
	endcase
end
endmodule

module layer1_N4_rsh_2(address, data);
input wire [5:0] address;
output reg [0:0] data;

always @(*) begin
	case(address)
		6'd0: data = 1'd0;
		6'd1: data = 1'd1;
		6'd2: data = 1'd1;
		6'd3: data = 1'd1;
		6'd4: data = 1'd0;
		6'd5: data = 1'd1;
		6'd6: data = 1'd1;
		6'd7: data = 1'd1;
		6'd8: data = 1'd0;
		6'd9: data = 1'd0;
		6'd10: data = 1'd1;
		6'd11: data = 1'd1;
		6'd12: data = 1'd0;
		6'd13: data = 1'd0;
		6'd14: data = 1'd1;
		6'd15: data = 1'd1;
		6'd16: data = 1'd0;
		6'd17: data = 1'd0;
		6'd18: data = 1'd1;
		6'd19: data = 1'd1;
		6'd20: data = 1'd0;
		6'd21: data = 1'd0;
		6'd22: data = 1'd1;
		6'd23: data = 1'd1;
		6'd24: data = 1'd0;
		6'd25: data = 1'd0;
		6'd26: data = 1'd1;
		6'd27: data = 1'd1;
		6'd28: data = 1'd0;
		6'd29: data = 1'd0;
		6'd30: data = 1'd0;
		6'd31: data = 1'd0;
		6'd32: data = 1'd1;
		6'd33: data = 1'd0;
		6'd34: data = 1'd0;
		6'd35: data = 1'd0;
		6'd36: data = 1'd1;
		6'd37: data = 1'd0;
		6'd38: data = 1'd0;
		6'd39: data = 1'd0;
		6'd40: data = 1'd1;
		6'd41: data = 1'd0;
		6'd42: data = 1'd0;
		6'd43: data = 1'd0;
		6'd44: data = 1'd1;
		6'd45: data = 1'd0;
		6'd46: data = 1'd0;
		6'd47: data = 1'd0;
		6'd48: data = 1'd1;
		6'd49: data = 1'd0;
		6'd50: data = 1'd0;
		6'd51: data = 1'd0;
		6'd52: data = 1'd1;
		6'd53: data = 1'd0;
		6'd54: data = 1'd0;
		6'd55: data = 1'd0;
		6'd56: data = 1'd1;
		6'd57: data = 1'd1;
		6'd58: data = 1'd0;
		6'd59: data = 1'd0;
		6'd60: data = 1'd1;
		6'd61: data = 1'd1;
		6'd62: data = 1'd0;
		6'd63: data = 1'd0;
		default: data = 1'd0;
	endcase
end
endmodule

module layer1_N4_lb_2(address, data);
input wire [9:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		10'd0: data = 3'd7;
		10'd1: data = 3'd6;
		10'd2: data = 3'd2;
		10'd3: data = 3'd7;
		10'd4: data = 3'd7;
		10'd5: data = 3'd4;
		10'd6: data = 3'd1;
		10'd7: data = 3'd6;
		10'd8: data = 3'd5;
		10'd9: data = 3'd2;
		10'd10: data = 3'd0;
		10'd11: data = 3'd5;
		10'd12: data = 3'd2;
		10'd13: data = 3'd0;
		10'd14: data = 3'd7;
		10'd15: data = 3'd4;
		10'd16: data = 3'd6;
		10'd17: data = 3'd5;
		10'd18: data = 3'd6;
		10'd19: data = 3'd3;
		10'd20: data = 3'd2;
		10'd21: data = 3'd1;
		10'd22: data = 3'd5;
		10'd23: data = 3'd2;
		10'd24: data = 3'd0;
		10'd25: data = 3'd0;
		10'd26: data = 3'd4;
		10'd27: data = 3'd1;
		10'd28: data = 3'd0;
		10'd29: data = 3'd0;
		10'd30: data = 3'd3;
		10'd31: data = 3'd0;
		10'd32: data = 3'd0;
		10'd33: data = 3'd0;
		10'd34: data = 3'd3;
		10'd35: data = 3'd0;
		10'd36: data = 3'd0;
		10'd37: data = 3'd0;
		10'd38: data = 3'd3;
		10'd39: data = 3'd0;
		10'd40: data = 3'd0;
		10'd41: data = 3'd0;
		10'd42: data = 3'd3;
		10'd43: data = 3'd0;
		10'd44: data = 3'd0;
		10'd45: data = 3'd0;
		10'd46: data = 3'd3;
		10'd47: data = 3'd0;
		10'd48: data = 3'd0;
		10'd49: data = 3'd0;
		10'd50: data = 3'd3;
		10'd51: data = 3'd0;
		10'd52: data = 3'd0;
		10'd53: data = 3'd0;
		10'd54: data = 3'd3;
		10'd55: data = 3'd0;
		10'd56: data = 3'd0;
		10'd57: data = 3'd0;
		10'd58: data = 3'd2;
		10'd59: data = 3'd0;
		10'd60: data = 3'd0;
		10'd61: data = 3'd0;
		10'd62: data = 3'd2;
		10'd63: data = 3'd1;
		10'd64: data = 3'd7;
		10'd65: data = 3'd6;
		10'd66: data = 3'd2;
		10'd67: data = 3'd7;
		10'd68: data = 3'd7;
		10'd69: data = 3'd4;
		10'd70: data = 3'd1;
		10'd71: data = 3'd6;
		10'd72: data = 3'd5;
		10'd73: data = 3'd2;
		10'd74: data = 3'd0;
		10'd75: data = 3'd6;
		10'd76: data = 3'd3;
		10'd77: data = 3'd0;
		10'd78: data = 3'd0;
		10'd79: data = 3'd5;
		10'd80: data = 3'd7;
		10'd81: data = 3'd6;
		10'd82: data = 3'd7;
		10'd83: data = 3'd4;
		10'd84: data = 3'd3;
		10'd85: data = 3'd2;
		10'd86: data = 3'd6;
		10'd87: data = 3'd2;
		10'd88: data = 3'd0;
		10'd89: data = 3'd0;
		10'd90: data = 3'd4;
		10'd91: data = 3'd1;
		10'd92: data = 3'd0;
		10'd93: data = 3'd0;
		10'd94: data = 3'd4;
		10'd95: data = 3'd0;
		10'd96: data = 3'd0;
		10'd97: data = 3'd0;
		10'd98: data = 3'd3;
		10'd99: data = 3'd0;
		10'd100: data = 3'd0;
		10'd101: data = 3'd0;
		10'd102: data = 3'd3;
		10'd103: data = 3'd0;
		10'd104: data = 3'd0;
		10'd105: data = 3'd0;
		10'd106: data = 3'd4;
		10'd107: data = 3'd0;
		10'd108: data = 3'd0;
		10'd109: data = 3'd0;
		10'd110: data = 3'd4;
		10'd111: data = 3'd0;
		10'd112: data = 3'd0;
		10'd113: data = 3'd0;
		10'd114: data = 3'd4;
		10'd115: data = 3'd0;
		10'd116: data = 3'd0;
		10'd117: data = 3'd1;
		10'd118: data = 3'd3;
		10'd119: data = 3'd0;
		10'd120: data = 3'd0;
		10'd121: data = 3'd1;
		10'd122: data = 3'd3;
		10'd123: data = 3'd1;
		10'd124: data = 3'd0;
		10'd125: data = 3'd1;
		10'd126: data = 3'd3;
		10'd127: data = 3'd2;
		10'd128: data = 3'd7;
		10'd129: data = 3'd6;
		10'd130: data = 3'd2;
		10'd131: data = 3'd0;
		10'd132: data = 3'd7;
		10'd133: data = 3'd4;
		10'd134: data = 3'd2;
		10'd135: data = 3'd7;
		10'd136: data = 3'd5;
		10'd137: data = 3'd2;
		10'd138: data = 3'd1;
		10'd139: data = 3'd6;
		10'd140: data = 3'd3;
		10'd141: data = 3'd1;
		10'd142: data = 3'd0;
		10'd143: data = 3'd5;
		10'd144: data = 3'd0;
		10'd145: data = 3'd7;
		10'd146: data = 3'd7;
		10'd147: data = 3'd4;
		10'd148: data = 3'd4;
		10'd149: data = 3'd3;
		10'd150: data = 3'd6;
		10'd151: data = 3'd3;
		10'd152: data = 3'd0;
		10'd153: data = 3'd0;
		10'd154: data = 3'd5;
		10'd155: data = 3'd1;
		10'd156: data = 3'd0;
		10'd157: data = 3'd0;
		10'd158: data = 3'd4;
		10'd159: data = 3'd0;
		10'd160: data = 3'd0;
		10'd161: data = 3'd1;
		10'd162: data = 3'd3;
		10'd163: data = 3'd0;
		10'd164: data = 3'd0;
		10'd165: data = 3'd1;
		10'd166: data = 3'd4;
		10'd167: data = 3'd0;
		10'd168: data = 3'd0;
		10'd169: data = 3'd1;
		10'd170: data = 3'd5;
		10'd171: data = 3'd0;
		10'd172: data = 3'd0;
		10'd173: data = 3'd1;
		10'd174: data = 3'd5;
		10'd175: data = 3'd0;
		10'd176: data = 3'd0;
		10'd177: data = 3'd2;
		10'd178: data = 3'd4;
		10'd179: data = 3'd0;
		10'd180: data = 3'd0;
		10'd181: data = 3'd2;
		10'd182: data = 3'd4;
		10'd183: data = 3'd1;
		10'd184: data = 3'd1;
		10'd185: data = 3'd2;
		10'd186: data = 3'd4;
		10'd187: data = 3'd1;
		10'd188: data = 3'd1;
		10'd189: data = 3'd2;
		10'd190: data = 3'd3;
		10'd191: data = 3'd2;
		10'd192: data = 3'd7;
		10'd193: data = 3'd6;
		10'd194: data = 3'd3;
		10'd195: data = 3'd1;
		10'd196: data = 3'd7;
		10'd197: data = 3'd4;
		10'd198: data = 3'd2;
		10'd199: data = 3'd0;
		10'd200: data = 3'd5;
		10'd201: data = 3'd3;
		10'd202: data = 3'd1;
		10'd203: data = 3'd7;
		10'd204: data = 3'd3;
		10'd205: data = 3'd1;
		10'd206: data = 3'd0;
		10'd207: data = 3'd6;
		10'd208: data = 3'd1;
		10'd209: data = 3'd0;
		10'd210: data = 3'd0;
		10'd211: data = 3'd4;
		10'd212: data = 3'd5;
		10'd213: data = 3'd5;
		10'd214: data = 3'd7;
		10'd215: data = 3'd3;
		10'd216: data = 3'd1;
		10'd217: data = 3'd2;
		10'd218: data = 3'd6;
		10'd219: data = 3'd2;
		10'd220: data = 3'd0;
		10'd221: data = 3'd1;
		10'd222: data = 3'd4;
		10'd223: data = 3'd0;
		10'd224: data = 3'd0;
		10'd225: data = 3'd1;
		10'd226: data = 3'd4;
		10'd227: data = 3'd0;
		10'd228: data = 3'd0;
		10'd229: data = 3'd2;
		10'd230: data = 3'd4;
		10'd231: data = 3'd0;
		10'd232: data = 3'd0;
		10'd233: data = 3'd2;
		10'd234: data = 3'd5;
		10'd235: data = 3'd0;
		10'd236: data = 3'd0;
		10'd237: data = 3'd2;
		10'd238: data = 3'd5;
		10'd239: data = 3'd0;
		10'd240: data = 3'd0;
		10'd241: data = 3'd3;
		10'd242: data = 3'd5;
		10'd243: data = 3'd1;
		10'd244: data = 3'd1;
		10'd245: data = 3'd3;
		10'd246: data = 3'd5;
		10'd247: data = 3'd1;
		10'd248: data = 3'd1;
		10'd249: data = 3'd3;
		10'd250: data = 3'd4;
		10'd251: data = 3'd2;
		10'd252: data = 3'd2;
		10'd253: data = 3'd3;
		10'd254: data = 3'd4;
		10'd255: data = 3'd3;
		10'd256: data = 3'd7;
		10'd257: data = 3'd7;
		10'd258: data = 3'd3;
		10'd259: data = 3'd1;
		10'd260: data = 3'd7;
		10'd261: data = 3'd5;
		10'd262: data = 3'd3;
		10'd263: data = 3'd0;
		10'd264: data = 3'd5;
		10'd265: data = 3'd3;
		10'd266: data = 3'd2;
		10'd267: data = 3'd0;
		10'd268: data = 3'd3;
		10'd269: data = 3'd2;
		10'd270: data = 3'd1;
		10'd271: data = 3'd6;
		10'd272: data = 3'd1;
		10'd273: data = 3'd0;
		10'd274: data = 3'd0;
		10'd275: data = 3'd5;
		10'd276: data = 3'd6;
		10'd277: data = 3'd6;
		10'd278: data = 3'd7;
		10'd279: data = 3'd3;
		10'd280: data = 3'd2;
		10'd281: data = 3'd3;
		10'd282: data = 3'd6;
		10'd283: data = 3'd2;
		10'd284: data = 3'd0;
		10'd285: data = 3'd2;
		10'd286: data = 3'd5;
		10'd287: data = 3'd1;
		10'd288: data = 3'd0;
		10'd289: data = 3'd2;
		10'd290: data = 3'd4;
		10'd291: data = 3'd0;
		10'd292: data = 3'd0;
		10'd293: data = 3'd2;
		10'd294: data = 3'd5;
		10'd295: data = 3'd0;
		10'd296: data = 3'd1;
		10'd297: data = 3'd3;
		10'd298: data = 3'd6;
		10'd299: data = 3'd0;
		10'd300: data = 3'd1;
		10'd301: data = 3'd3;
		10'd302: data = 3'd6;
		10'd303: data = 3'd0;
		10'd304: data = 3'd1;
		10'd305: data = 3'd3;
		10'd306: data = 3'd6;
		10'd307: data = 3'd1;
		10'd308: data = 3'd1;
		10'd309: data = 3'd4;
		10'd310: data = 3'd6;
		10'd311: data = 3'd2;
		10'd312: data = 3'd2;
		10'd313: data = 3'd4;
		10'd314: data = 3'd5;
		10'd315: data = 3'd2;
		10'd316: data = 3'd2;
		10'd317: data = 3'd4;
		10'd318: data = 3'd5;
		10'd319: data = 3'd3;
		10'd320: data = 3'd7;
		10'd321: data = 3'd7;
		10'd322: data = 3'd4;
		10'd323: data = 3'd2;
		10'd324: data = 3'd7;
		10'd325: data = 3'd6;
		10'd326: data = 3'd3;
		10'd327: data = 3'd1;
		10'd328: data = 3'd5;
		10'd329: data = 3'd4;
		10'd330: data = 3'd2;
		10'd331: data = 3'd0;
		10'd332: data = 3'd3;
		10'd333: data = 3'd2;
		10'd334: data = 3'd1;
		10'd335: data = 3'd7;
		10'd336: data = 3'd1;
		10'd337: data = 3'd1;
		10'd338: data = 3'd1;
		10'd339: data = 3'd5;
		10'd340: data = 3'd7;
		10'd341: data = 3'd7;
		10'd342: data = 3'd0;
		10'd343: data = 3'd4;
		10'd344: data = 3'd4;
		10'd345: data = 3'd5;
		10'd346: data = 3'd6;
		10'd347: data = 3'd2;
		10'd348: data = 3'd1;
		10'd349: data = 3'd3;
		10'd350: data = 3'd5;
		10'd351: data = 3'd1;
		10'd352: data = 3'd1;
		10'd353: data = 3'd3;
		10'd354: data = 3'd5;
		10'd355: data = 3'd0;
		10'd356: data = 3'd1;
		10'd357: data = 3'd3;
		10'd358: data = 3'd5;
		10'd359: data = 3'd0;
		10'd360: data = 3'd1;
		10'd361: data = 3'd3;
		10'd362: data = 3'd6;
		10'd363: data = 3'd0;
		10'd364: data = 3'd1;
		10'd365: data = 3'd4;
		10'd366: data = 3'd7;
		10'd367: data = 3'd1;
		10'd368: data = 3'd2;
		10'd369: data = 3'd4;
		10'd370: data = 3'd7;
		10'd371: data = 3'd2;
		10'd372: data = 3'd2;
		10'd373: data = 3'd4;
		10'd374: data = 3'd6;
		10'd375: data = 3'd2;
		10'd376: data = 3'd2;
		10'd377: data = 3'd5;
		10'd378: data = 3'd6;
		10'd379: data = 3'd3;
		10'd380: data = 3'd3;
		10'd381: data = 3'd5;
		10'd382: data = 3'd6;
		10'd383: data = 3'd4;
		10'd384: data = 3'd7;
		10'd385: data = 3'd7;
		10'd386: data = 3'd4;
		10'd387: data = 3'd3;
		10'd388: data = 3'd7;
		10'd389: data = 3'd6;
		10'd390: data = 3'd3;
		10'd391: data = 3'd2;
		10'd392: data = 3'd6;
		10'd393: data = 3'd4;
		10'd394: data = 3'd3;
		10'd395: data = 3'd0;
		10'd396: data = 3'd3;
		10'd397: data = 3'd3;
		10'd398: data = 3'd2;
		10'd399: data = 3'd7;
		10'd400: data = 3'd1;
		10'd401: data = 3'd1;
		10'd402: data = 3'd1;
		10'd403: data = 3'd6;
		10'd404: data = 3'd7;
		10'd405: data = 3'd0;
		10'd406: data = 3'd0;
		10'd407: data = 3'd4;
		10'd408: data = 3'd5;
		10'd409: data = 3'd7;
		10'd410: data = 3'd7;
		10'd411: data = 3'd3;
		10'd412: data = 3'd2;
		10'd413: data = 3'd5;
		10'd414: data = 3'd6;
		10'd415: data = 3'd1;
		10'd416: data = 3'd1;
		10'd417: data = 3'd4;
		10'd418: data = 3'd6;
		10'd419: data = 3'd0;
		10'd420: data = 3'd1;
		10'd421: data = 3'd4;
		10'd422: data = 3'd6;
		10'd423: data = 3'd0;
		10'd424: data = 3'd1;
		10'd425: data = 3'd4;
		10'd426: data = 3'd7;
		10'd427: data = 3'd1;
		10'd428: data = 3'd2;
		10'd429: data = 3'd4;
		10'd430: data = 3'd7;
		10'd431: data = 3'd1;
		10'd432: data = 3'd2;
		10'd433: data = 3'd5;
		10'd434: data = 3'd7;
		10'd435: data = 3'd2;
		10'd436: data = 3'd3;
		10'd437: data = 3'd5;
		10'd438: data = 3'd7;
		10'd439: data = 3'd3;
		10'd440: data = 3'd3;
		10'd441: data = 3'd5;
		10'd442: data = 3'd7;
		10'd443: data = 3'd3;
		10'd444: data = 3'd3;
		10'd445: data = 3'd6;
		10'd446: data = 3'd7;
		10'd447: data = 3'd4;
		10'd448: data = 3'd7;
		10'd449: data = 3'd7;
		10'd450: data = 3'd5;
		10'd451: data = 3'd3;
		10'd452: data = 3'd7;
		10'd453: data = 3'd6;
		10'd454: data = 3'd4;
		10'd455: data = 3'd2;
		10'd456: data = 3'd6;
		10'd457: data = 3'd5;
		10'd458: data = 3'd3;
		10'd459: data = 3'd1;
		10'd460: data = 3'd3;
		10'd461: data = 3'd3;
		10'd462: data = 3'd2;
		10'd463: data = 3'd7;
		10'd464: data = 3'd1;
		10'd465: data = 3'd2;
		10'd466: data = 3'd1;
		10'd467: data = 3'd6;
		10'd468: data = 3'd0;
		10'd469: data = 3'd1;
		10'd470: data = 3'd0;
		10'd471: data = 3'd5;
		10'd472: data = 3'd6;
		10'd473: data = 3'd0;
		10'd474: data = 3'd7;
		10'd475: data = 3'd3;
		10'd476: data = 3'd3;
		10'd477: data = 3'd6;
		10'd478: data = 3'd7;
		10'd479: data = 3'd2;
		10'd480: data = 3'd2;
		10'd481: data = 3'd5;
		10'd482: data = 3'd7;
		10'd483: data = 3'd1;
		10'd484: data = 3'd1;
		10'd485: data = 3'd5;
		10'd486: data = 3'd7;
		10'd487: data = 3'd1;
		10'd488: data = 3'd2;
		10'd489: data = 3'd5;
		10'd490: data = 3'd7;
		10'd491: data = 3'd1;
		10'd492: data = 3'd2;
		10'd493: data = 3'd5;
		10'd494: data = 3'd0;
		10'd495: data = 3'd2;
		10'd496: data = 3'd3;
		10'd497: data = 3'd5;
		10'd498: data = 3'd0;
		10'd499: data = 3'd3;
		10'd500: data = 3'd3;
		10'd501: data = 3'd5;
		10'd502: data = 3'd0;
		10'd503: data = 3'd3;
		10'd504: data = 3'd3;
		10'd505: data = 3'd6;
		10'd506: data = 3'd0;
		10'd507: data = 3'd4;
		10'd508: data = 3'd4;
		10'd509: data = 3'd6;
		10'd510: data = 3'd0;
		10'd511: data = 3'd5;
		10'd512: data = 3'd7;
		10'd513: data = 3'd7;
		10'd514: data = 3'd5;
		10'd515: data = 3'd4;
		10'd516: data = 3'd7;
		10'd517: data = 3'd7;
		10'd518: data = 3'd4;
		10'd519: data = 3'd3;
		10'd520: data = 3'd6;
		10'd521: data = 3'd5;
		10'd522: data = 3'd3;
		10'd523: data = 3'd1;
		10'd524: data = 3'd3;
		10'd525: data = 3'd4;
		10'd526: data = 3'd3;
		10'd527: data = 3'd0;
		10'd528: data = 3'd2;
		10'd529: data = 3'd3;
		10'd530: data = 3'd1;
		10'd531: data = 3'd6;
		10'd532: data = 3'd0;
		10'd533: data = 3'd2;
		10'd534: data = 3'd1;
		10'd535: data = 3'd5;
		10'd536: data = 3'd7;
		10'd537: data = 3'd1;
		10'd538: data = 3'd0;
		10'd539: data = 3'd4;
		10'd540: data = 3'd4;
		10'd541: data = 3'd7;
		10'd542: data = 3'd0;
		10'd543: data = 3'd2;
		10'd544: data = 3'd2;
		10'd545: data = 3'd7;
		10'd546: data = 3'd0;
		10'd547: data = 3'd2;
		10'd548: data = 3'd2;
		10'd549: data = 3'd6;
		10'd550: data = 3'd7;
		10'd551: data = 3'd2;
		10'd552: data = 3'd2;
		10'd553: data = 3'd6;
		10'd554: data = 3'd0;
		10'd555: data = 3'd2;
		10'd556: data = 3'd3;
		10'd557: data = 3'd5;
		10'd558: data = 3'd0;
		10'd559: data = 3'd2;
		10'd560: data = 3'd3;
		10'd561: data = 3'd5;
		10'd562: data = 3'd0;
		10'd563: data = 3'd3;
		10'd564: data = 3'd4;
		10'd565: data = 3'd6;
		10'd566: data = 3'd0;
		10'd567: data = 3'd4;
		10'd568: data = 3'd4;
		10'd569: data = 3'd6;
		10'd570: data = 3'd0;
		10'd571: data = 3'd4;
		10'd572: data = 3'd4;
		10'd573: data = 3'd6;
		10'd574: data = 3'd0;
		10'd575: data = 3'd5;
		10'd576: data = 3'd7;
		10'd577: data = 3'd7;
		10'd578: data = 3'd5;
		10'd579: data = 3'd4;
		10'd580: data = 3'd7;
		10'd581: data = 3'd7;
		10'd582: data = 3'd5;
		10'd583: data = 3'd3;
		10'd584: data = 3'd5;
		10'd585: data = 3'd6;
		10'd586: data = 3'd4;
		10'd587: data = 3'd2;
		10'd588: data = 3'd4;
		10'd589: data = 3'd4;
		10'd590: data = 3'd3;
		10'd591: data = 3'd0;
		10'd592: data = 3'd2;
		10'd593: data = 3'd3;
		10'd594: data = 3'd2;
		10'd595: data = 3'd7;
		10'd596: data = 3'd1;
		10'd597: data = 3'd3;
		10'd598: data = 3'd1;
		10'd599: data = 3'd5;
		10'd600: data = 3'd7;
		10'd601: data = 3'd2;
		10'd602: data = 3'd1;
		10'd603: data = 3'd4;
		10'd604: data = 3'd5;
		10'd605: data = 3'd1;
		10'd606: data = 3'd1;
		10'd607: data = 3'd3;
		10'd608: data = 3'd3;
		10'd609: data = 3'd0;
		10'd610: data = 3'd0;
		10'd611: data = 3'd3;
		10'd612: data = 3'd3;
		10'd613: data = 3'd0;
		10'd614: data = 3'd0;
		10'd615: data = 3'd3;
		10'd616: data = 3'd3;
		10'd617: data = 3'd6;
		10'd618: data = 3'd0;
		10'd619: data = 3'd2;
		10'd620: data = 3'd3;
		10'd621: data = 3'd6;
		10'd622: data = 3'd0;
		10'd623: data = 3'd3;
		10'd624: data = 3'd4;
		10'd625: data = 3'd6;
		10'd626: data = 3'd0;
		10'd627: data = 3'd4;
		10'd628: data = 3'd4;
		10'd629: data = 3'd6;
		10'd630: data = 3'd0;
		10'd631: data = 3'd4;
		10'd632: data = 3'd4;
		10'd633: data = 3'd6;
		10'd634: data = 3'd0;
		10'd635: data = 3'd5;
		10'd636: data = 3'd4;
		10'd637: data = 3'd6;
		10'd638: data = 3'd0;
		10'd639: data = 3'd5;
		10'd640: data = 3'd7;
		10'd641: data = 3'd7;
		10'd642: data = 3'd6;
		10'd643: data = 3'd4;
		10'd644: data = 3'd6;
		10'd645: data = 3'd7;
		10'd646: data = 3'd5;
		10'd647: data = 3'd3;
		10'd648: data = 3'd5;
		10'd649: data = 3'd6;
		10'd650: data = 3'd4;
		10'd651: data = 3'd2;
		10'd652: data = 3'd4;
		10'd653: data = 3'd5;
		10'd654: data = 3'd3;
		10'd655: data = 3'd0;
		10'd656: data = 3'd2;
		10'd657: data = 3'd4;
		10'd658: data = 3'd2;
		10'd659: data = 3'd7;
		10'd660: data = 3'd1;
		10'd661: data = 3'd3;
		10'd662: data = 3'd2;
		10'd663: data = 3'd6;
		10'd664: data = 3'd0;
		10'd665: data = 3'd3;
		10'd666: data = 3'd2;
		10'd667: data = 3'd5;
		10'd668: data = 3'd6;
		10'd669: data = 3'd2;
		10'd670: data = 3'd2;
		10'd671: data = 3'd4;
		10'd672: data = 3'd5;
		10'd673: data = 3'd2;
		10'd674: data = 3'd1;
		10'd675: data = 3'd4;
		10'd676: data = 3'd4;
		10'd677: data = 3'd1;
		10'd678: data = 3'd1;
		10'd679: data = 3'd3;
		10'd680: data = 3'd4;
		10'd681: data = 3'd7;
		10'd682: data = 3'd1;
		10'd683: data = 3'd3;
		10'd684: data = 3'd4;
		10'd685: data = 3'd6;
		10'd686: data = 3'd1;
		10'd687: data = 3'd3;
		10'd688: data = 3'd4;
		10'd689: data = 3'd6;
		10'd690: data = 3'd0;
		10'd691: data = 3'd4;
		10'd692: data = 3'd4;
		10'd693: data = 3'd6;
		10'd694: data = 3'd0;
		10'd695: data = 3'd4;
		10'd696: data = 3'd5;
		10'd697: data = 3'd6;
		10'd698: data = 3'd0;
		10'd699: data = 3'd5;
		10'd700: data = 3'd5;
		10'd701: data = 3'd6;
		10'd702: data = 3'd0;
		10'd703: data = 3'd5;
		10'd704: data = 3'd7;
		10'd705: data = 3'd7;
		10'd706: data = 3'd6;
		10'd707: data = 3'd4;
		10'd708: data = 3'd6;
		10'd709: data = 3'd7;
		10'd710: data = 3'd5;
		10'd711: data = 3'd3;
		10'd712: data = 3'd5;
		10'd713: data = 3'd7;
		10'd714: data = 3'd4;
		10'd715: data = 3'd2;
		10'd716: data = 3'd4;
		10'd717: data = 3'd6;
		10'd718: data = 3'd4;
		10'd719: data = 3'd1;
		10'd720: data = 3'd3;
		10'd721: data = 3'd5;
		10'd722: data = 3'd3;
		10'd723: data = 3'd7;
		10'd724: data = 3'd1;
		10'd725: data = 3'd4;
		10'd726: data = 3'd3;
		10'd727: data = 3'd6;
		10'd728: data = 3'd0;
		10'd729: data = 3'd3;
		10'd730: data = 3'd3;
		10'd731: data = 3'd6;
		10'd732: data = 3'd7;
		10'd733: data = 3'd3;
		10'd734: data = 3'd2;
		10'd735: data = 3'd5;
		10'd736: data = 3'd6;
		10'd737: data = 3'd3;
		10'd738: data = 3'd2;
		10'd739: data = 3'd5;
		10'd740: data = 3'd5;
		10'd741: data = 3'd1;
		10'd742: data = 3'd1;
		10'd743: data = 3'd4;
		10'd744: data = 3'd5;
		10'd745: data = 3'd0;
		10'd746: data = 3'd1;
		10'd747: data = 3'd4;
		10'd748: data = 3'd5;
		10'd749: data = 3'd7;
		10'd750: data = 3'd1;
		10'd751: data = 3'd4;
		10'd752: data = 3'd5;
		10'd753: data = 3'd7;
		10'd754: data = 3'd1;
		10'd755: data = 3'd4;
		10'd756: data = 3'd5;
		10'd757: data = 3'd6;
		10'd758: data = 3'd0;
		10'd759: data = 3'd4;
		10'd760: data = 3'd5;
		10'd761: data = 3'd6;
		10'd762: data = 3'd0;
		10'd763: data = 3'd5;
		10'd764: data = 3'd5;
		10'd765: data = 3'd6;
		10'd766: data = 3'd0;
		10'd767: data = 3'd6;
		10'd768: data = 3'd6;
		10'd769: data = 3'd7;
		10'd770: data = 3'd7;
		10'd771: data = 3'd4;
		10'd772: data = 3'd5;
		10'd773: data = 3'd7;
		10'd774: data = 3'd6;
		10'd775: data = 3'd3;
		10'd776: data = 3'd4;
		10'd777: data = 3'd7;
		10'd778: data = 3'd5;
		10'd779: data = 3'd2;
		10'd780: data = 3'd4;
		10'd781: data = 3'd6;
		10'd782: data = 3'd4;
		10'd783: data = 3'd1;
		10'd784: data = 3'd3;
		10'd785: data = 3'd6;
		10'd786: data = 3'd4;
		10'd787: data = 3'd7;
		10'd788: data = 3'd2;
		10'd789: data = 3'd5;
		10'd790: data = 3'd4;
		10'd791: data = 3'd7;
		10'd792: data = 3'd1;
		10'd793: data = 3'd4;
		10'd794: data = 3'd3;
		10'd795: data = 3'd6;
		10'd796: data = 3'd0;
		10'd797: data = 3'd4;
		10'd798: data = 3'd3;
		10'd799: data = 3'd6;
		10'd800: data = 3'd0;
		10'd801: data = 3'd3;
		10'd802: data = 3'd3;
		10'd803: data = 3'd5;
		10'd804: data = 3'd7;
		10'd805: data = 3'd2;
		10'd806: data = 3'd2;
		10'd807: data = 3'd5;
		10'd808: data = 3'd7;
		10'd809: data = 3'd1;
		10'd810: data = 3'd2;
		10'd811: data = 3'd4;
		10'd812: data = 3'd6;
		10'd813: data = 3'd0;
		10'd814: data = 3'd2;
		10'd815: data = 3'd4;
		10'd816: data = 3'd6;
		10'd817: data = 3'd7;
		10'd818: data = 3'd2;
		10'd819: data = 3'd4;
		10'd820: data = 3'd6;
		10'd821: data = 3'd7;
		10'd822: data = 3'd1;
		10'd823: data = 3'd4;
		10'd824: data = 3'd6;
		10'd825: data = 3'd7;
		10'd826: data = 3'd0;
		10'd827: data = 3'd5;
		10'd828: data = 3'd6;
		10'd829: data = 3'd7;
		10'd830: data = 3'd0;
		10'd831: data = 3'd6;
		10'd832: data = 3'd6;
		10'd833: data = 3'd7;
		10'd834: data = 3'd7;
		10'd835: data = 3'd4;
		10'd836: data = 3'd5;
		10'd837: data = 3'd7;
		10'd838: data = 3'd6;
		10'd839: data = 3'd3;
		10'd840: data = 3'd4;
		10'd841: data = 3'd7;
		10'd842: data = 3'd5;
		10'd843: data = 3'd2;
		10'd844: data = 3'd3;
		10'd845: data = 3'd7;
		10'd846: data = 3'd5;
		10'd847: data = 3'd1;
		10'd848: data = 3'd3;
		10'd849: data = 3'd6;
		10'd850: data = 3'd5;
		10'd851: data = 3'd0;
		10'd852: data = 3'd2;
		10'd853: data = 3'd6;
		10'd854: data = 3'd5;
		10'd855: data = 3'd0;
		10'd856: data = 3'd2;
		10'd857: data = 3'd5;
		10'd858: data = 3'd4;
		10'd859: data = 3'd7;
		10'd860: data = 3'd1;
		10'd861: data = 3'd5;
		10'd862: data = 3'd4;
		10'd863: data = 3'd7;
		10'd864: data = 3'd1;
		10'd865: data = 3'd4;
		10'd866: data = 3'd4;
		10'd867: data = 3'd6;
		10'd868: data = 3'd1;
		10'd869: data = 3'd3;
		10'd870: data = 3'd3;
		10'd871: data = 3'd6;
		10'd872: data = 3'd0;
		10'd873: data = 3'd2;
		10'd874: data = 3'd3;
		10'd875: data = 3'd5;
		10'd876: data = 3'd0;
		10'd877: data = 3'd1;
		10'd878: data = 3'd3;
		10'd879: data = 3'd5;
		10'd880: data = 3'd0;
		10'd881: data = 3'd0;
		10'd882: data = 3'd2;
		10'd883: data = 3'd5;
		10'd884: data = 3'd0;
		10'd885: data = 3'd0;
		10'd886: data = 3'd1;
		10'd887: data = 3'd5;
		10'd888: data = 3'd0;
		10'd889: data = 3'd0;
		10'd890: data = 3'd1;
		10'd891: data = 3'd5;
		10'd892: data = 3'd0;
		10'd893: data = 3'd0;
		10'd894: data = 3'd1;
		10'd895: data = 3'd6;
		10'd896: data = 3'd5;
		10'd897: data = 3'd7;
		10'd898: data = 3'd7;
		10'd899: data = 3'd5;
		10'd900: data = 3'd4;
		10'd901: data = 3'd7;
		10'd902: data = 3'd7;
		10'd903: data = 3'd3;
		10'd904: data = 3'd3;
		10'd905: data = 3'd7;
		10'd906: data = 3'd6;
		10'd907: data = 3'd2;
		10'd908: data = 3'd3;
		10'd909: data = 3'd7;
		10'd910: data = 3'd6;
		10'd911: data = 3'd2;
		10'd912: data = 3'd3;
		10'd913: data = 3'd7;
		10'd914: data = 3'd6;
		10'd915: data = 3'd1;
		10'd916: data = 3'd3;
		10'd917: data = 3'd6;
		10'd918: data = 3'd5;
		10'd919: data = 3'd1;
		10'd920: data = 3'd3;
		10'd921: data = 3'd6;
		10'd922: data = 3'd5;
		10'd923: data = 3'd0;
		10'd924: data = 3'd3;
		10'd925: data = 3'd5;
		10'd926: data = 3'd5;
		10'd927: data = 3'd0;
		10'd928: data = 3'd3;
		10'd929: data = 3'd5;
		10'd930: data = 3'd4;
		10'd931: data = 3'd7;
		10'd932: data = 3'd3;
		10'd933: data = 3'd5;
		10'd934: data = 3'd4;
		10'd935: data = 3'd7;
		10'd936: data = 3'd2;
		10'd937: data = 3'd4;
		10'd938: data = 3'd3;
		10'd939: data = 3'd6;
		10'd940: data = 3'd2;
		10'd941: data = 3'd3;
		10'd942: data = 3'd3;
		10'd943: data = 3'd6;
		10'd944: data = 3'd2;
		10'd945: data = 3'd2;
		10'd946: data = 3'd3;
		10'd947: data = 3'd6;
		10'd948: data = 3'd1;
		10'd949: data = 3'd1;
		10'd950: data = 3'd2;
		10'd951: data = 3'd5;
		10'd952: data = 3'd1;
		10'd953: data = 3'd1;
		10'd954: data = 3'd1;
		10'd955: data = 3'd5;
		10'd956: data = 3'd1;
		10'd957: data = 3'd1;
		10'd958: data = 3'd1;
		10'd959: data = 3'd6;
		10'd960: data = 3'd5;
		10'd961: data = 3'd7;
		10'd962: data = 3'd7;
		10'd963: data = 3'd5;
		10'd964: data = 3'd4;
		10'd965: data = 3'd7;
		10'd966: data = 3'd7;
		10'd967: data = 3'd4;
		10'd968: data = 3'd3;
		10'd969: data = 3'd7;
		10'd970: data = 3'd7;
		10'd971: data = 3'd3;
		10'd972: data = 3'd3;
		10'd973: data = 3'd7;
		10'd974: data = 3'd7;
		10'd975: data = 3'd2;
		10'd976: data = 3'd3;
		10'd977: data = 3'd7;
		10'd978: data = 3'd7;
		10'd979: data = 3'd2;
		10'd980: data = 3'd4;
		10'd981: data = 3'd7;
		10'd982: data = 3'd6;
		10'd983: data = 3'd1;
		10'd984: data = 3'd4;
		10'd985: data = 3'd7;
		10'd986: data = 3'd6;
		10'd987: data = 3'd1;
		10'd988: data = 3'd4;
		10'd989: data = 3'd6;
		10'd990: data = 3'd6;
		10'd991: data = 3'd0;
		10'd992: data = 3'd5;
		10'd993: data = 3'd6;
		10'd994: data = 3'd5;
		10'd995: data = 3'd0;
		10'd996: data = 3'd5;
		10'd997: data = 3'd6;
		10'd998: data = 3'd5;
		10'd999: data = 3'd7;
		10'd1000: data = 3'd4;
		10'd1001: data = 3'd5;
		10'd1002: data = 3'd4;
		10'd1003: data = 3'd7;
		10'd1004: data = 3'd4;
		10'd1005: data = 3'd4;
		10'd1006: data = 3'd4;
		10'd1007: data = 3'd6;
		10'd1008: data = 3'd3;
		10'd1009: data = 3'd3;
		10'd1010: data = 3'd4;
		10'd1011: data = 3'd6;
		10'd1012: data = 3'd3;
		10'd1013: data = 3'd3;
		10'd1014: data = 3'd3;
		10'd1015: data = 3'd6;
		10'd1016: data = 3'd2;
		10'd1017: data = 3'd2;
		10'd1018: data = 3'd3;
		10'd1019: data = 3'd6;
		10'd1020: data = 3'd2;
		10'd1021: data = 3'd2;
		10'd1022: data = 3'd2;
		10'd1023: data = 3'd6;
		default: data = 3'd0;
	endcase
end
endmodule

module layer1_N4_2(address, data);
input wire [9:0] address;
output reg [3:0] data;

wire [4:0] i; layer1_N4_idx_2 idx_2_inst(address[9:4], i);
wire [0:0] t; layer1_N4_rsh_2 rsh_2_inst(address[9:4], t);
wire [0:0] b; layer1_N4_3 layer1_N4_3_inst(address[9:4], b);
wire [2:0] lb; layer1_N4_lb_2 lb_2_inst(address, lb);
wire [0:0] u; layer1_N4_ust_2 ust_2_inst({i, address[3:0]}, u);

always @(*) begin
	data = {(u >> t) + b, lb};
end
endmodule

module layer1_N4_ust_1(address, data);
input wire [7:0] address;
output reg [2:0] data;

always @(*) begin
	case(address)
		8'd0: data = 3'd3;
		8'd1: data = 3'd2;
		8'd2: data = 3'd1;
		8'd3: data = 3'd0;
		8'd4: data = 3'd0;
		8'd5: data = 3'd1;
		8'd6: data = 3'd2;
		8'd7: data = 3'd3;
		8'd8: data = 3'd4;
		8'd9: data = 3'd3;
		8'd10: data = 3'd2;
		8'd11: data = 3'd0;
		8'd12: data = 3'd0;
		8'd13: data = 3'd1;
		8'd14: data = 3'd2;
		8'd15: data = 3'd4;
		8'd16: data = 3'd4;
		8'd17: data = 3'd3;
		8'd18: data = 3'd1;
		8'd19: data = 3'd0;
		8'd20: data = 3'd2;
		8'd21: data = 3'd2;
		8'd22: data = 3'd1;
		8'd23: data = 3'd0;
		8'd24: data = 3'd0;
		8'd25: data = 3'd1;
		8'd26: data = 3'd2;
		8'd27: data = 3'd2;
		8'd28: data = 3'd0;
		8'd29: data = 3'd2;
		8'd30: data = 3'd3;
		8'd31: data = 3'd4;
		8'd32: data = 3'd4;
		8'd33: data = 3'd2;
		8'd34: data = 3'd1;
		8'd35: data = 3'd0;
		8'd36: data = 3'd0;
		8'd37: data = 3'd2;
		8'd38: data = 3'd2;
		8'd39: data = 3'd3;
		8'd40: data = 3'd2;
		8'd41: data = 3'd3;
		8'd42: data = 3'd2;
		8'd43: data = 3'd0;
		8'd44: data = 3'd1;
		8'd45: data = 3'd2;
		8'd46: data = 3'd2;
		8'd47: data = 3'd0;
		8'd48: data = 3'd0;
		8'd49: data = 3'd1;
		8'd50: data = 3'd2;
		8'd51: data = 3'd1;
		8'd52: data = 3'd5;
		8'd53: data = 3'd3;
		8'd54: data = 3'd2;
		8'd55: data = 3'd0;
		8'd56: data = 3'd2;
		8'd57: data = 3'd1;
		8'd58: data = 3'd0;
		8'd59: data = 3'd2;
		8'd60: data = 3'd0;
		8'd61: data = 3'd0;
		8'd62: data = 3'd1;
		8'd63: data = 3'd3;
		8'd64: data = 3'd1;
		8'd65: data = 3'd2;
		8'd66: data = 3'd1;
		8'd67: data = 3'd0;
		8'd68: data = 3'd2;
		8'd69: data = 3'd1;
		8'd70: data = 3'd0;
		8'd71: data = 3'd1;
		8'd72: data = 3'd0;
		8'd73: data = 3'd1;
		8'd74: data = 3'd1;
		8'd75: data = 3'd3;
		8'd76: data = 3'd1;
		8'd77: data = 3'd0;
		8'd78: data = 3'd1;
		8'd79: data = 3'd2;
		8'd80: data = 3'd0;
		8'd81: data = 3'd0;
		8'd82: data = 3'd1;
		8'd83: data = 3'd4;
		8'd84: data = 3'd1;
		8'd85: data = 3'd0;
		8'd86: data = 3'd1;
		8'd87: data = 3'd1;
		8'd88: data = 3'd0;
		8'd89: data = 3'd1;
		8'd90: data = 3'd3;
		8'd91: data = 3'd4;
		8'd92: data = 3'd3;
		8'd93: data = 3'd3;
		8'd94: data = 3'd2;
		8'd95: data = 3'd0;
		8'd96: data = 3'd0;
		8'd97: data = 3'd1;
		8'd98: data = 3'd2;
		8'd99: data = 3'd0;
		8'd100: data = 3'd2;
		8'd101: data = 3'd3;
		8'd102: data = 3'd1;
		8'd103: data = 3'd0;
		8'd104: data = 3'd1;
		8'd105: data = 3'd1;
		8'd106: data = 3'd0;
		8'd107: data = 3'd1;
		8'd108: data = 3'd3;
		8'd109: data = 3'd3;
		8'd110: data = 3'd1;
		8'd111: data = 3'd0;
		8'd112: data = 3'd3;
		8'd113: data = 3'd2;
		8'd114: data = 3'd0;
		8'd115: data = 3'd0;
		8'd116: data = 3'd1;
		8'd117: data = 3'd0;
		8'd118: data = 3'd0;
		8'd119: data = 3'd2;
		8'd120: data = 3'd0;
		8'd121: data = 3'd0;
		8'd122: data = 3'd2;
		8'd123: data = 3'd5;
		8'd124: data = 3'd3;
		8'd125: data = 3'd1;
		8'd126: data = 3'd0;
		8'd127: data = 3'd0;
		8'd128: data = 3'd0;
		8'd129: data = 3'd1;
		8'd130: data = 3'd2;
		8'd131: data = 3'd5;
		8'd132: data = 3'd0;
		8'd133: data = 3'd2;
		8'd134: data = 3'd2;
		8'd135: data = 3'd0;
		8'd136: data = 3'd3;
		8'd137: data = 3'd2;
		8'd138: data = 3'd2;
		8'd139: data = 3'd0;
		8'd140: data = 3'd2;
		8'd141: data = 3'd2;
		8'd142: data = 3'd2;
		8'd143: data = 3'd0;
		8'd144: data = 3'd0;
		8'd145: data = 3'd0;
		8'd146: data = 3'd2;
		8'd147: data = 3'd3;
		8'd148: data = 3'd0;
		8'd149: data = 3'd1;
		8'd150: data = 3'd0;
		8'd151: data = 3'd1;
		8'd152: data = 3'd3;
		8'd153: data = 3'd1;
		8'd154: data = 3'd1;
		8'd155: data = 3'd0;
		8'd156: data = 3'd1;
		8'd157: data = 3'd3;
		8'd158: data = 3'd2;
		8'd159: data = 3'd0;
		8'd160: data = 3'd1;
		8'd161: data = 3'd3;
		8'd162: data = 3'd1;
		8'd163: data = 3'd0;
		8'd164: data = 3'd0;
		8'd165: data = 3'd0;
		8'd166: data = 3'd2;
		8'd167: data = 3'd2;
		8'd168: data = 3'd2;
		8'd169: data = 3'd0;
		8'd170: data = 3'd0;
		8'd171: data = 3'd0;
		default: data = 3'd0;
	endcase
end
endmodule

module layer1_N4_idx_1(address, data);
input wire [9:0] address;
output reg [5:0] data;

always @(*) begin
	case(address)
		10'd0: data = 6'd0;
		10'd1: data = 6'd0;
		10'd2: data = 6'd2;
		10'd3: data = 6'd4;
		10'd4: data = 6'd0;
		10'd5: data = 6'd17;
		10'd6: data = 6'd0;
		10'd7: data = 6'd4;
		10'd8: data = 6'd5;
		10'd9: data = 6'd17;
		10'd10: data = 6'd0;
		10'd11: data = 6'd4;
		10'd12: data = 6'd5;
		10'd13: data = 6'd29;
		10'd14: data = 6'd0;
		10'd15: data = 6'd2;
		10'd16: data = 6'd5;
		10'd17: data = 6'd15;
		10'd18: data = 6'd0;
		10'd19: data = 6'd2;
		10'd20: data = 6'd0;
		10'd21: data = 6'd30;
		10'd22: data = 6'd0;
		10'd23: data = 6'd2;
		10'd24: data = 6'd2;
		10'd25: data = 6'd15;
		10'd26: data = 6'd5;
		10'd27: data = 6'd5;
		10'd28: data = 6'd0;
		10'd29: data = 6'd3;
		10'd30: data = 6'd11;
		10'd31: data = 6'd0;
		10'd32: data = 6'd0;
		10'd33: data = 6'd3;
		10'd34: data = 6'd11;
		10'd35: data = 6'd2;
		10'd36: data = 6'd0;
		10'd37: data = 6'd3;
		10'd38: data = 6'd11;
		10'd39: data = 6'd4;
		10'd40: data = 6'd0;
		10'd41: data = 6'd3;
		10'd42: data = 6'd12;
		10'd43: data = 6'd4;
		10'd44: data = 6'd0;
		10'd45: data = 6'd3;
		10'd46: data = 6'd12;
		10'd47: data = 6'd31;
		10'd48: data = 6'd0;
		10'd49: data = 6'd3;
		10'd50: data = 6'd6;
		10'd51: data = 6'd0;
		10'd52: data = 6'd0;
		10'd53: data = 6'd20;
		10'd54: data = 6'd3;
		10'd55: data = 6'd4;
		10'd56: data = 6'd0;
		10'd57: data = 6'd3;
		10'd58: data = 6'd1;
		10'd59: data = 6'd13;
		10'd60: data = 6'd0;
		10'd61: data = 6'd3;
		10'd62: data = 6'd1;
		10'd63: data = 6'd2;
		10'd64: data = 6'd0;
		10'd65: data = 6'd0;
		10'd66: data = 6'd0;
		10'd67: data = 6'd2;
		10'd68: data = 6'd0;
		10'd69: data = 6'd17;
		10'd70: data = 6'd0;
		10'd71: data = 6'd2;
		10'd72: data = 6'd5;
		10'd73: data = 6'd14;
		10'd74: data = 6'd0;
		10'd75: data = 6'd0;
		10'd76: data = 6'd5;
		10'd77: data = 6'd14;
		10'd78: data = 6'd2;
		10'd79: data = 6'd4;
		10'd80: data = 6'd5;
		10'd81: data = 6'd15;
		10'd82: data = 6'd0;
		10'd83: data = 6'd2;
		10'd84: data = 6'd2;
		10'd85: data = 6'd30;
		10'd86: data = 6'd2;
		10'd87: data = 6'd0;
		10'd88: data = 6'd4;
		10'd89: data = 6'd20;
		10'd90: data = 6'd0;
		10'd91: data = 6'd0;
		10'd92: data = 6'd0;
		10'd93: data = 6'd3;
		10'd94: data = 6'd16;
		10'd95: data = 6'd0;
		10'd96: data = 6'd0;
		10'd97: data = 6'd3;
		10'd98: data = 6'd16;
		10'd99: data = 6'd2;
		10'd100: data = 6'd0;
		10'd101: data = 6'd3;
		10'd102: data = 6'd11;
		10'd103: data = 6'd4;
		10'd104: data = 6'd0;
		10'd105: data = 6'd3;
		10'd106: data = 6'd24;
		10'd107: data = 6'd31;
		10'd108: data = 6'd0;
		10'd109: data = 6'd18;
		10'd110: data = 6'd12;
		10'd111: data = 6'd28;
		10'd112: data = 6'd0;
		10'd113: data = 6'd18;
		10'd114: data = 6'd1;
		10'd115: data = 6'd4;
		10'd116: data = 6'd0;
		10'd117: data = 6'd3;
		10'd118: data = 6'd1;
		10'd119: data = 6'd13;
		10'd120: data = 6'd3;
		10'd121: data = 6'd3;
		10'd122: data = 6'd1;
		10'd123: data = 6'd4;
		10'd124: data = 6'd3;
		10'd125: data = 6'd3;
		10'd126: data = 6'd7;
		10'd127: data = 6'd4;
		10'd128: data = 6'd0;
		10'd129: data = 6'd0;
		10'd130: data = 6'd0;
		10'd131: data = 6'd4;
		10'd132: data = 6'd0;
		10'd133: data = 6'd17;
		10'd134: data = 6'd0;
		10'd135: data = 6'd2;
		10'd136: data = 6'd5;
		10'd137: data = 6'd14;
		10'd138: data = 6'd0;
		10'd139: data = 6'd2;
		10'd140: data = 6'd5;
		10'd141: data = 6'd29;
		10'd142: data = 6'd0;
		10'd143: data = 6'd2;
		10'd144: data = 6'd2;
		10'd145: data = 6'd15;
		10'd146: data = 6'd0;
		10'd147: data = 6'd5;
		10'd148: data = 6'd2;
		10'd149: data = 6'd32;
		10'd150: data = 6'd0;
		10'd151: data = 6'd2;
		10'd152: data = 6'd0;
		10'd153: data = 6'd32;
		10'd154: data = 6'd0;
		10'd155: data = 6'd0;
		10'd156: data = 6'd0;
		10'd157: data = 6'd1;
		10'd158: data = 6'd16;
		10'd159: data = 6'd0;
		10'd160: data = 6'd0;
		10'd161: data = 6'd3;
		10'd162: data = 6'd10;
		10'd163: data = 6'd2;
		10'd164: data = 6'd0;
		10'd165: data = 6'd18;
		10'd166: data = 6'd16;
		10'd167: data = 6'd4;
		10'd168: data = 6'd3;
		10'd169: data = 6'd18;
		10'd170: data = 6'd11;
		10'd171: data = 6'd28;
		10'd172: data = 6'd1;
		10'd173: data = 6'd18;
		10'd174: data = 6'd11;
		10'd175: data = 6'd8;
		10'd176: data = 6'd1;
		10'd177: data = 6'd1;
		10'd178: data = 6'd6;
		10'd179: data = 6'd2;
		10'd180: data = 6'd9;
		10'd181: data = 6'd1;
		10'd182: data = 6'd1;
		10'd183: data = 6'd4;
		10'd184: data = 6'd3;
		10'd185: data = 6'd3;
		10'd186: data = 6'd6;
		10'd187: data = 6'd13;
		10'd188: data = 6'd1;
		10'd189: data = 6'd3;
		10'd190: data = 6'd1;
		10'd191: data = 6'd2;
		10'd192: data = 6'd0;
		10'd193: data = 6'd0;
		10'd194: data = 6'd0;
		10'd195: data = 6'd2;
		10'd196: data = 6'd0;
		10'd197: data = 6'd17;
		10'd198: data = 6'd0;
		10'd199: data = 6'd0;
		10'd200: data = 6'd5;
		10'd201: data = 6'd14;
		10'd202: data = 6'd0;
		10'd203: data = 6'd0;
		10'd204: data = 6'd5;
		10'd205: data = 6'd19;
		10'd206: data = 6'd0;
		10'd207: data = 6'd2;
		10'd208: data = 6'd2;
		10'd209: data = 6'd20;
		10'd210: data = 6'd0;
		10'd211: data = 6'd0;
		10'd212: data = 6'd2;
		10'd213: data = 6'd3;
		10'd214: data = 6'd0;
		10'd215: data = 6'd0;
		10'd216: data = 6'd0;
		10'd217: data = 6'd3;
		10'd218: data = 6'd2;
		10'd219: data = 6'd2;
		10'd220: data = 6'd2;
		10'd221: data = 6'd3;
		10'd222: data = 6'd5;
		10'd223: data = 6'd0;
		10'd224: data = 6'd3;
		10'd225: data = 6'd3;
		10'd226: data = 6'd25;
		10'd227: data = 6'd2;
		10'd228: data = 6'd3;
		10'd229: data = 6'd18;
		10'd230: data = 6'd10;
		10'd231: data = 6'd28;
		10'd232: data = 6'd1;
		10'd233: data = 6'd1;
		10'd234: data = 6'd11;
		10'd235: data = 6'd8;
		10'd236: data = 6'd7;
		10'd237: data = 6'd6;
		10'd238: data = 6'd12;
		10'd239: data = 6'd4;
		10'd240: data = 6'd6;
		10'd241: data = 6'd1;
		10'd242: data = 6'd12;
		10'd243: data = 6'd4;
		10'd244: data = 6'd3;
		10'd245: data = 6'd1;
		10'd246: data = 6'd6;
		10'd247: data = 6'd13;
		10'd248: data = 6'd7;
		10'd249: data = 6'd1;
		10'd250: data = 6'd1;
		10'd251: data = 6'd4;
		10'd252: data = 6'd1;
		10'd253: data = 6'd37;
		10'd254: data = 6'd1;
		10'd255: data = 6'd4;
		10'd256: data = 6'd0;
		10'd257: data = 6'd0;
		10'd258: data = 6'd0;
		10'd259: data = 6'd2;
		10'd260: data = 6'd0;
		10'd261: data = 6'd14;
		10'd262: data = 6'd2;
		10'd263: data = 6'd2;
		10'd264: data = 6'd5;
		10'd265: data = 6'd21;
		10'd266: data = 6'd5;
		10'd267: data = 6'd0;
		10'd268: data = 6'd5;
		10'd269: data = 6'd3;
		10'd270: data = 6'd0;
		10'd271: data = 6'd5;
		10'd272: data = 6'd0;
		10'd273: data = 6'd7;
		10'd274: data = 6'd0;
		10'd275: data = 6'd5;
		10'd276: data = 6'd2;
		10'd277: data = 6'd1;
		10'd278: data = 6'd0;
		10'd279: data = 6'd0;
		10'd280: data = 6'd0;
		10'd281: data = 6'd22;
		10'd282: data = 6'd0;
		10'd283: data = 6'd0;
		10'd284: data = 6'd26;
		10'd285: data = 6'd22;
		10'd286: data = 6'd0;
		10'd287: data = 6'd2;
		10'd288: data = 6'd21;
		10'd289: data = 6'd3;
		10'd290: data = 6'd23;
		10'd291: data = 6'd38;
		10'd292: data = 6'd19;
		10'd293: data = 6'd3;
		10'd294: data = 6'd25;
		10'd295: data = 6'd0;
		10'd296: data = 6'd3;
		10'd297: data = 6'd1;
		10'd298: data = 6'd11;
		10'd299: data = 6'd4;
		10'd300: data = 6'd1;
		10'd301: data = 6'd6;
		10'd302: data = 6'd24;
		10'd303: data = 6'd13;
		10'd304: data = 6'd7;
		10'd305: data = 6'd6;
		10'd306: data = 6'd12;
		10'd307: data = 6'd2;
		10'd308: data = 6'd6;
		10'd309: data = 6'd1;
		10'd310: data = 6'd3;
		10'd311: data = 6'd4;
		10'd312: data = 6'd3;
		10'd313: data = 6'd1;
		10'd314: data = 6'd1;
		10'd315: data = 6'd13;
		10'd316: data = 6'd6;
		10'd317: data = 6'd9;
		10'd318: data = 6'd1;
		10'd319: data = 6'd2;
		10'd320: data = 6'd0;
		10'd321: data = 6'd0;
		10'd322: data = 6'd5;
		10'd323: data = 6'd0;
		10'd324: data = 6'd0;
		10'd325: data = 6'd2;
		10'd326: data = 6'd0;
		10'd327: data = 6'd2;
		10'd328: data = 6'd5;
		10'd329: data = 6'd3;
		10'd330: data = 6'd0;
		10'd331: data = 6'd2;
		10'd332: data = 6'd5;
		10'd333: data = 6'd7;
		10'd334: data = 6'd0;
		10'd335: data = 6'd4;
		10'd336: data = 6'd0;
		10'd337: data = 6'd3;
		10'd338: data = 6'd2;
		10'd339: data = 6'd0;
		10'd340: data = 6'd4;
		10'd341: data = 6'd1;
		10'd342: data = 6'd0;
		10'd343: data = 6'd5;
		10'd344: data = 6'd2;
		10'd345: data = 6'd1;
		10'd346: data = 6'd2;
		10'd347: data = 6'd0;
		10'd348: data = 6'd14;
		10'd349: data = 6'd7;
		10'd350: data = 6'd2;
		10'd351: data = 6'd0;
		10'd352: data = 6'd3;
		10'd353: data = 6'd3;
		10'd354: data = 6'd27;
		10'd355: data = 6'd0;
		10'd356: data = 6'd1;
		10'd357: data = 6'd1;
		10'd358: data = 6'd10;
		10'd359: data = 6'd4;
		10'd360: data = 6'd3;
		10'd361: data = 6'd1;
		10'd362: data = 6'd11;
		10'd363: data = 6'd13;
		10'd364: data = 6'd7;
		10'd365: data = 6'd7;
		10'd366: data = 6'd11;
		10'd367: data = 6'd4;
		10'd368: data = 6'd1;
		10'd369: data = 6'd7;
		10'd370: data = 6'd12;
		10'd371: data = 6'd4;
		10'd372: data = 6'd7;
		10'd373: data = 6'd6;
		10'd374: data = 6'd6;
		10'd375: data = 6'd13;
		10'd376: data = 6'd6;
		10'd377: data = 6'd1;
		10'd378: data = 6'd1;
		10'd379: data = 6'd4;
		10'd380: data = 6'd3;
		10'd381: data = 6'd9;
		10'd382: data = 6'd7;
		10'd383: data = 6'd4;
		10'd384: data = 6'd0;
		10'd385: data = 6'd0;
		10'd386: data = 6'd0;
		10'd387: data = 6'd0;
		10'd388: data = 6'd0;
		10'd389: data = 6'd14;
		10'd390: data = 6'd0;
		10'd391: data = 6'd0;
		10'd392: data = 6'd10;
		10'd393: data = 6'd19;
		10'd394: data = 6'd4;
		10'd395: data = 6'd5;
		10'd396: data = 6'd5;
		10'd397: data = 6'd3;
		10'd398: data = 6'd5;
		10'd399: data = 6'd0;
		10'd400: data = 6'd0;
		10'd401: data = 6'd1;
		10'd402: data = 6'd0;
		10'd403: data = 6'd4;
		10'd404: data = 6'd0;
		10'd405: data = 6'd1;
		10'd406: data = 6'd0;
		10'd407: data = 6'd0;
		10'd408: data = 6'd14;
		10'd409: data = 6'd1;
		10'd410: data = 6'd8;
		10'd411: data = 6'd0;
		10'd412: data = 6'd14;
		10'd413: data = 6'd3;
		10'd414: data = 6'd4;
		10'd415: data = 6'd8;
		10'd416: data = 6'd3;
		10'd417: data = 6'd22;
		10'd418: data = 6'd27;
		10'd419: data = 6'd4;
		10'd420: data = 6'd3;
		10'd421: data = 6'd1;
		10'd422: data = 6'd25;
		10'd423: data = 6'd2;
		10'd424: data = 6'd7;
		10'd425: data = 6'd1;
		10'd426: data = 6'd16;
		10'd427: data = 6'd4;
		10'd428: data = 6'd3;
		10'd429: data = 6'd1;
		10'd430: data = 6'd11;
		10'd431: data = 6'd13;
		10'd432: data = 6'd7;
		10'd433: data = 6'd3;
		10'd434: data = 6'd12;
		10'd435: data = 6'd2;
		10'd436: data = 6'd1;
		10'd437: data = 6'd3;
		10'd438: data = 6'd6;
		10'd439: data = 6'd4;
		10'd440: data = 6'd7;
		10'd441: data = 6'd7;
		10'd442: data = 6'd6;
		10'd443: data = 6'd13;
		10'd444: data = 6'd6;
		10'd445: data = 6'd1;
		10'd446: data = 6'd3;
		10'd447: data = 6'd2;
		10'd448: data = 6'd0;
		10'd449: data = 6'd0;
		10'd450: data = 6'd4;
		10'd451: data = 6'd10;
		10'd452: data = 6'd0;
		10'd453: data = 6'd21;
		10'd454: data = 6'd5;
		10'd455: data = 6'd10;
		10'd456: data = 6'd10;
		10'd457: data = 6'd1;
		10'd458: data = 6'd0;
		10'd459: data = 6'd5;
		10'd460: data = 6'd5;
		10'd461: data = 6'd1;
		10'd462: data = 6'd0;
		10'd463: data = 6'd0;
		10'd464: data = 6'd0;
		10'd465: data = 6'd6;
		10'd466: data = 6'd0;
		10'd467: data = 6'd0;
		10'd468: data = 6'd4;
		10'd469: data = 6'd1;
		10'd470: data = 6'd4;
		10'd471: data = 6'd4;
		10'd472: data = 6'd14;
		10'd473: data = 6'd1;
		10'd474: data = 6'd2;
		10'd475: data = 6'd0;
		10'd476: data = 6'd19;
		10'd477: data = 6'd22;
		10'd478: data = 6'd8;
		10'd479: data = 6'd0;
		10'd480: data = 6'd3;
		10'd481: data = 6'd7;
		10'd482: data = 6'd0;
		10'd483: data = 6'd4;
		10'd484: data = 6'd1;
		10'd485: data = 6'd1;
		10'd486: data = 6'd5;
		10'd487: data = 6'd4;
		10'd488: data = 6'd3;
		10'd489: data = 6'd6;
		10'd490: data = 6'd39;
		10'd491: data = 6'd13;
		10'd492: data = 6'd7;
		10'd493: data = 6'd7;
		10'd494: data = 6'd11;
		10'd495: data = 6'd4;
		10'd496: data = 6'd1;
		10'd497: data = 6'd7;
		10'd498: data = 6'd24;
		10'd499: data = 6'd4;
		10'd500: data = 6'd7;
		10'd501: data = 6'd7;
		10'd502: data = 6'd12;
		10'd503: data = 6'd13;
		10'd504: data = 6'd6;
		10'd505: data = 6'd1;
		10'd506: data = 6'd3;
		10'd507: data = 6'd4;
		10'd508: data = 6'd1;
		10'd509: data = 6'd1;
		10'd510: data = 6'd3;
		10'd511: data = 6'd4;
		10'd512: data = 6'd0;
		10'd513: data = 6'd0;
		10'd514: data = 6'd5;
		10'd515: data = 6'd0;
		10'd516: data = 6'd0;
		10'd517: data = 6'd0;
		10'd518: data = 6'd0;
		10'd519: data = 6'd0;
		10'd520: data = 6'd0;
		10'd521: data = 6'd6;
		10'd522: data = 6'd0;
		10'd523: data = 6'd5;
		10'd524: data = 6'd5;
		10'd525: data = 6'd7;
		10'd526: data = 6'd4;
		10'd527: data = 6'd2;
		10'd528: data = 6'd0;
		10'd529: data = 6'd3;
		10'd530: data = 6'd2;
		10'd531: data = 6'd0;
		10'd532: data = 6'd17;
		10'd533: data = 6'd1;
		10'd534: data = 6'd0;
		10'd535: data = 6'd0;
		10'd536: data = 6'd14;
		10'd537: data = 6'd1;
		10'd538: data = 6'd4;
		10'd539: data = 6'd0;
		10'd540: data = 6'd3;
		10'd541: data = 6'd7;
		10'd542: data = 6'd0;
		10'd543: data = 6'd2;
		10'd544: data = 6'd3;
		10'd545: data = 6'd1;
		10'd546: data = 6'd5;
		10'd547: data = 6'd4;
		10'd548: data = 6'd1;
		10'd549: data = 6'd1;
		10'd550: data = 6'd10;
		10'd551: data = 6'd4;
		10'd552: data = 6'd1;
		10'd553: data = 6'd3;
		10'd554: data = 6'd16;
		10'd555: data = 6'd4;
		10'd556: data = 6'd3;
		10'd557: data = 6'd6;
		10'd558: data = 6'd33;
		10'd559: data = 6'd13;
		10'd560: data = 6'd7;
		10'd561: data = 6'd6;
		10'd562: data = 6'd12;
		10'd563: data = 6'd2;
		10'd564: data = 6'd1;
		10'd565: data = 6'd1;
		10'd566: data = 6'd12;
		10'd567: data = 6'd4;
		10'd568: data = 6'd1;
		10'd569: data = 6'd1;
		10'd570: data = 6'd3;
		10'd571: data = 6'd13;
		10'd572: data = 6'd1;
		10'd573: data = 6'd1;
		10'd574: data = 6'd3;
		10'd575: data = 6'd2;
		10'd576: data = 6'd0;
		10'd577: data = 6'd0;
		10'd578: data = 6'd5;
		10'd579: data = 6'd0;
		10'd580: data = 6'd0;
		10'd581: data = 6'd0;
		10'd582: data = 6'd4;
		10'd583: data = 6'd0;
		10'd584: data = 6'd10;
		10'd585: data = 6'd1;
		10'd586: data = 6'd5;
		10'd587: data = 6'd0;
		10'd588: data = 6'd0;
		10'd589: data = 6'd6;
		10'd590: data = 6'd0;
		10'd591: data = 6'd5;
		10'd592: data = 6'd0;
		10'd593: data = 6'd1;
		10'd594: data = 6'd0;
		10'd595: data = 6'd2;
		10'd596: data = 6'd14;
		10'd597: data = 6'd7;
		10'd598: data = 6'd4;
		10'd599: data = 6'd0;
		10'd600: data = 6'd19;
		10'd601: data = 6'd6;
		10'd602: data = 6'd0;
		10'd603: data = 6'd4;
		10'd604: data = 6'd15;
		10'd605: data = 6'd6;
		10'd606: data = 6'd0;
		10'd607: data = 6'd2;
		10'd608: data = 6'd7;
		10'd609: data = 6'd1;
		10'd610: data = 6'd23;
		10'd611: data = 6'd4;
		10'd612: data = 6'd1;
		10'd613: data = 6'd3;
		10'd614: data = 6'd10;
		10'd615: data = 6'd8;
		10'd616: data = 6'd1;
		10'd617: data = 6'd6;
		10'd618: data = 6'd40;
		10'd619: data = 6'd13;
		10'd620: data = 6'd6;
		10'd621: data = 6'd3;
		10'd622: data = 6'd33;
		10'd623: data = 6'd4;
		10'd624: data = 6'd1;
		10'd625: data = 6'd3;
		10'd626: data = 6'd12;
		10'd627: data = 6'd8;
		10'd628: data = 6'd1;
		10'd629: data = 6'd1;
		10'd630: data = 6'd12;
		10'd631: data = 6'd2;
		10'd632: data = 6'd9;
		10'd633: data = 6'd1;
		10'd634: data = 6'd6;
		10'd635: data = 6'd8;
		10'd636: data = 6'd9;
		10'd637: data = 6'd1;
		10'd638: data = 6'd3;
		10'd639: data = 6'd2;
		10'd640: data = 6'd0;
		10'd641: data = 6'd0;
		10'd642: data = 6'd10;
		10'd643: data = 6'd10;
		10'd644: data = 6'd0;
		10'd645: data = 6'd0;
		10'd646: data = 6'd5;
		10'd647: data = 6'd4;
		10'd648: data = 6'd0;
		10'd649: data = 6'd9;
		10'd650: data = 6'd0;
		10'd651: data = 6'd0;
		10'd652: data = 6'd0;
		10'd653: data = 6'd6;
		10'd654: data = 6'd27;
		10'd655: data = 6'd5;
		10'd656: data = 6'd26;
		10'd657: data = 6'd6;
		10'd658: data = 6'd2;
		10'd659: data = 6'd2;
		10'd660: data = 6'd21;
		10'd661: data = 6'd1;
		10'd662: data = 6'd0;
		10'd663: data = 6'd0;
		10'd664: data = 6'd3;
		10'd665: data = 6'd7;
		10'd666: data = 6'd0;
		10'd667: data = 6'd8;
		10'd668: data = 6'd1;
		10'd669: data = 6'd6;
		10'd670: data = 6'd5;
		10'd671: data = 6'd2;
		10'd672: data = 6'd1;
		10'd673: data = 6'd3;
		10'd674: data = 6'd0;
		10'd675: data = 6'd8;
		10'd676: data = 6'd3;
		10'd677: data = 6'd1;
		10'd678: data = 6'd5;
		10'd679: data = 6'd2;
		10'd680: data = 6'd1;
		10'd681: data = 6'd6;
		10'd682: data = 6'd16;
		10'd683: data = 6'd2;
		10'd684: data = 6'd7;
		10'd685: data = 6'd6;
		10'd686: data = 6'd11;
		10'd687: data = 6'd4;
		10'd688: data = 6'd7;
		10'd689: data = 6'd7;
		10'd690: data = 6'd12;
		10'd691: data = 6'd8;
		10'd692: data = 6'd7;
		10'd693: data = 6'd9;
		10'd694: data = 6'd6;
		10'd695: data = 6'd2;
		10'd696: data = 6'd3;
		10'd697: data = 6'd9;
		10'd698: data = 6'd6;
		10'd699: data = 6'd4;
		10'd700: data = 6'd3;
		10'd701: data = 6'd9;
		10'd702: data = 6'd3;
		10'd703: data = 6'd2;
		10'd704: data = 6'd0;
		10'd705: data = 6'd0;
		10'd706: data = 6'd10;
		10'd707: data = 6'd2;
		10'd708: data = 6'd0;
		10'd709: data = 6'd0;
		10'd710: data = 6'd5;
		10'd711: data = 6'd2;
		10'd712: data = 6'd3;
		10'd713: data = 6'd0;
		10'd714: data = 6'd0;
		10'd715: data = 6'd4;
		10'd716: data = 6'd3;
		10'd717: data = 6'd9;
		10'd718: data = 6'd0;
		10'd719: data = 6'd0;
		10'd720: data = 6'd3;
		10'd721: data = 6'd6;
		10'd722: data = 6'd0;
		10'd723: data = 6'd0;
		10'd724: data = 6'd19;
		10'd725: data = 6'd1;
		10'd726: data = 6'd0;
		10'd727: data = 6'd4;
		10'd728: data = 6'd6;
		10'd729: data = 6'd1;
		10'd730: data = 6'd5;
		10'd731: data = 6'd8;
		10'd732: data = 6'd1;
		10'd733: data = 6'd7;
		10'd734: data = 6'd27;
		10'd735: data = 6'd4;
		10'd736: data = 6'd3;
		10'd737: data = 6'd1;
		10'd738: data = 6'd0;
		10'd739: data = 6'd8;
		10'd740: data = 6'd7;
		10'd741: data = 6'd6;
		10'd742: data = 6'd23;
		10'd743: data = 6'd4;
		10'd744: data = 6'd1;
		10'd745: data = 6'd6;
		10'd746: data = 6'd10;
		10'd747: data = 6'd4;
		10'd748: data = 6'd7;
		10'd749: data = 6'd6;
		10'd750: data = 6'd11;
		10'd751: data = 6'd8;
		10'd752: data = 6'd1;
		10'd753: data = 6'd1;
		10'd754: data = 6'd11;
		10'd755: data = 6'd8;
		10'd756: data = 6'd3;
		10'd757: data = 6'd7;
		10'd758: data = 6'd6;
		10'd759: data = 6'd2;
		10'd760: data = 6'd14;
		10'd761: data = 6'd7;
		10'd762: data = 6'd6;
		10'd763: data = 6'd4;
		10'd764: data = 6'd26;
		10'd765: data = 6'd7;
		10'd766: data = 6'd15;
		10'd767: data = 6'd8;
		10'd768: data = 6'd0;
		10'd769: data = 6'd0;
		10'd770: data = 6'd0;
		10'd771: data = 6'd2;
		10'd772: data = 6'd3;
		10'd773: data = 6'd0;
		10'd774: data = 6'd10;
		10'd775: data = 6'd2;
		10'd776: data = 6'd3;
		10'd777: data = 6'd0;
		10'd778: data = 6'd5;
		10'd779: data = 6'd2;
		10'd780: data = 6'd3;
		10'd781: data = 6'd9;
		10'd782: data = 6'd0;
		10'd783: data = 6'd4;
		10'd784: data = 6'd3;
		10'd785: data = 6'd9;
		10'd786: data = 6'd0;
		10'd787: data = 6'd2;
		10'd788: data = 6'd3;
		10'd789: data = 6'd6;
		10'd790: data = 6'd5;
		10'd791: data = 6'd4;
		10'd792: data = 6'd7;
		10'd793: data = 6'd6;
		10'd794: data = 6'd34;
		10'd795: data = 6'd2;
		10'd796: data = 6'd1;
		10'd797: data = 6'd7;
		10'd798: data = 6'd0;
		10'd799: data = 6'd4;
		10'd800: data = 6'd1;
		10'd801: data = 6'd6;
		10'd802: data = 6'd0;
		10'd803: data = 6'd2;
		10'd804: data = 6'd1;
		10'd805: data = 6'd6;
		10'd806: data = 6'd23;
		10'd807: data = 6'd4;
		10'd808: data = 6'd7;
		10'd809: data = 6'd6;
		10'd810: data = 6'd25;
		10'd811: data = 6'd13;
		10'd812: data = 6'd7;
		10'd813: data = 6'd7;
		10'd814: data = 6'd16;
		10'd815: data = 6'd2;
		10'd816: data = 6'd9;
		10'd817: data = 6'd7;
		10'd818: data = 6'd12;
		10'd819: data = 6'd2;
		10'd820: data = 6'd21;
		10'd821: data = 6'd1;
		10'd822: data = 6'd1;
		10'd823: data = 6'd2;
		10'd824: data = 6'd26;
		10'd825: data = 6'd3;
		10'd826: data = 6'd6;
		10'd827: data = 6'd4;
		10'd828: data = 6'd0;
		10'd829: data = 6'd3;
		10'd830: data = 6'd1;
		10'd831: data = 6'd8;
		10'd832: data = 6'd0;
		10'd833: data = 6'd0;
		10'd834: data = 6'd0;
		10'd835: data = 6'd5;
		10'd836: data = 6'd3;
		10'd837: data = 6'd0;
		10'd838: data = 6'd10;
		10'd839: data = 6'd2;
		10'd840: data = 6'd3;
		10'd841: data = 6'd0;
		10'd842: data = 6'd35;
		10'd843: data = 6'd2;
		10'd844: data = 6'd15;
		10'd845: data = 6'd0;
		10'd846: data = 6'd5;
		10'd847: data = 6'd0;
		10'd848: data = 6'd41;
		10'd849: data = 6'd9;
		10'd850: data = 6'd2;
		10'd851: data = 6'd2;
		10'd852: data = 6'd1;
		10'd853: data = 6'd9;
		10'd854: data = 6'd2;
		10'd855: data = 6'd0;
		10'd856: data = 6'd7;
		10'd857: data = 6'd7;
		10'd858: data = 6'd5;
		10'd859: data = 6'd2;
		10'd860: data = 6'd1;
		10'd861: data = 6'd1;
		10'd862: data = 6'd5;
		10'd863: data = 6'd8;
		10'd864: data = 6'd9;
		10'd865: data = 6'd7;
		10'd866: data = 6'd5;
		10'd867: data = 6'd2;
		10'd868: data = 6'd6;
		10'd869: data = 6'd6;
		10'd870: data = 6'd0;
		10'd871: data = 6'd8;
		10'd872: data = 6'd6;
		10'd873: data = 6'd7;
		10'd874: data = 6'd5;
		10'd875: data = 6'd2;
		10'd876: data = 6'd9;
		10'd877: data = 6'd7;
		10'd878: data = 6'd10;
		10'd879: data = 6'd4;
		10'd880: data = 6'd0;
		10'd881: data = 6'd7;
		10'd882: data = 6'd24;
		10'd883: data = 6'd4;
		10'd884: data = 6'd0;
		10'd885: data = 6'd3;
		10'd886: data = 6'd12;
		10'd887: data = 6'd8;
		10'd888: data = 6'd2;
		10'd889: data = 6'd0;
		10'd890: data = 6'd1;
		10'd891: data = 6'd4;
		10'd892: data = 6'd2;
		10'd893: data = 6'd0;
		10'd894: data = 6'd3;
		10'd895: data = 6'd8;
		10'd896: data = 6'd3;
		10'd897: data = 6'd0;
		10'd898: data = 6'd0;
		10'd899: data = 6'd0;
		10'd900: data = 6'd20;
		10'd901: data = 6'd0;
		10'd902: data = 6'd0;
		10'd903: data = 6'd5;
		10'd904: data = 6'd15;
		10'd905: data = 6'd0;
		10'd906: data = 6'd10;
		10'd907: data = 6'd0;
		10'd908: data = 6'd36;
		10'd909: data = 6'd0;
		10'd910: data = 6'd10;
		10'd911: data = 6'd0;
		10'd912: data = 6'd1;
		10'd913: data = 6'd0;
		10'd914: data = 6'd10;
		10'd915: data = 6'd4;
		10'd916: data = 6'd1;
		10'd917: data = 6'd9;
		10'd918: data = 6'd35;
		10'd919: data = 6'd0;
		10'd920: data = 6'd7;
		10'd921: data = 6'd9;
		10'd922: data = 6'd5;
		10'd923: data = 6'd4;
		10'd924: data = 6'd6;
		10'd925: data = 6'd6;
		10'd926: data = 6'd5;
		10'd927: data = 6'd8;
		10'd928: data = 6'd6;
		10'd929: data = 6'd3;
		10'd930: data = 6'd34;
		10'd931: data = 6'd4;
		10'd932: data = 6'd9;
		10'd933: data = 6'd3;
		10'd934: data = 6'd5;
		10'd935: data = 6'd8;
		10'd936: data = 6'd9;
		10'd937: data = 6'd3;
		10'd938: data = 6'd23;
		10'd939: data = 6'd4;
		10'd940: data = 6'd0;
		10'd941: data = 6'd3;
		10'd942: data = 6'd11;
		10'd943: data = 6'd8;
		10'd944: data = 6'd0;
		10'd945: data = 6'd3;
		10'd946: data = 6'd11;
		10'd947: data = 6'd8;
		10'd948: data = 6'd2;
		10'd949: data = 6'd1;
		10'd950: data = 6'd12;
		10'd951: data = 6'd13;
		10'd952: data = 6'd2;
		10'd953: data = 6'd0;
		10'd954: data = 6'd6;
		10'd955: data = 6'd2;
		10'd956: data = 6'd2;
		10'd957: data = 6'd0;
		10'd958: data = 6'd3;
		10'd959: data = 6'd8;
		10'd960: data = 6'd3;
		10'd961: data = 6'd0;
		10'd962: data = 6'd0;
		10'd963: data = 6'd4;
		10'd964: data = 6'd20;
		10'd965: data = 6'd0;
		10'd966: data = 6'd0;
		10'd967: data = 6'd4;
		10'd968: data = 6'd15;
		10'd969: data = 6'd0;
		10'd970: data = 6'd0;
		10'd971: data = 6'd0;
		10'd972: data = 6'd36;
		10'd973: data = 6'd0;
		10'd974: data = 6'd0;
		10'd975: data = 6'd2;
		10'd976: data = 6'd22;
		10'd977: data = 6'd0;
		10'd978: data = 6'd0;
		10'd979: data = 6'd0;
		10'd980: data = 6'd1;
		10'd981: data = 6'd0;
		10'd982: data = 6'd10;
		10'd983: data = 6'd2;
		10'd984: data = 6'd1;
		10'd985: data = 6'd0;
		10'd986: data = 6'd10;
		10'd987: data = 6'd4;
		10'd988: data = 6'd6;
		10'd989: data = 6'd9;
		10'd990: data = 6'd10;
		10'd991: data = 6'd2;
		10'd992: data = 6'd9;
		10'd993: data = 6'd1;
		10'd994: data = 6'd5;
		10'd995: data = 6'd4;
		10'd996: data = 6'd1;
		10'd997: data = 6'd3;
		10'd998: data = 6'd2;
		10'd999: data = 6'd2;
		10'd1000: data = 6'd1;
		10'd1001: data = 6'd1;
		10'd1002: data = 6'd5;
		10'd1003: data = 6'd4;
		10'd1004: data = 6'd0;
		10'd1005: data = 6'd1;
		10'd1006: data = 6'd16;
		10'd1007: data = 6'd2;
		10'd1008: data = 6'd0;
		10'd1009: data = 6'd9;
		10'd1010: data = 6'd11;
		10'd1011: data = 6'd2;
		10'd1012: data = 6'd0;
		10'd1013: data = 6'd0;
		10'd1014: data = 6'd9;
		10'd1015: data = 6'd4;
		10'd1016: data = 6'd2;
		10'd1017: data = 6'd3;
		10'd1018: data = 6'd0;
		10'd1019: data = 6'd4;
		10'd1020: data = 6'd42;
		10'd1021: data = 6'd0;
		10'd1022: data = 6'd3;
		10'd1023: data = 6'd4;
		default: data = 6'd0;
	endcase
end
endmodule

module layer1_N4_rsh_1(address, data);
input wire [9:0] address;
output reg [1:0] data;

always @(*) begin
	case(address)
		10'd0: data = 2'd2;
		10'd1: data = 2'd1;
		10'd2: data = 2'd1;
		10'd3: data = 2'd1;
		10'd4: data = 2'd2;
		10'd5: data = 2'd0;
		10'd6: data = 2'd0;
		10'd7: data = 2'd1;
		10'd8: data = 2'd0;
		10'd9: data = 2'd0;
		10'd10: data = 2'd0;
		10'd11: data = 2'd1;
		10'd12: data = 2'd0;
		10'd13: data = 2'd0;
		10'd14: data = 2'd0;
		10'd15: data = 2'd1;
		10'd16: data = 2'd0;
		10'd17: data = 2'd0;
		10'd18: data = 2'd0;
		10'd19: data = 2'd1;
		10'd20: data = 2'd0;
		10'd21: data = 2'd0;
		10'd22: data = 2'd0;
		10'd23: data = 2'd1;
		10'd24: data = 2'd2;
		10'd25: data = 2'd0;
		10'd26: data = 2'd0;
		10'd27: data = 2'd0;
		10'd28: data = 2'd2;
		10'd29: data = 2'd2;
		10'd30: data = 2'd1;
		10'd31: data = 2'd0;
		10'd32: data = 2'd2;
		10'd33: data = 2'd2;
		10'd34: data = 2'd1;
		10'd35: data = 2'd1;
		10'd36: data = 2'd2;
		10'd37: data = 2'd2;
		10'd38: data = 2'd1;
		10'd39: data = 2'd1;
		10'd40: data = 2'd2;
		10'd41: data = 2'd2;
		10'd42: data = 2'd0;
		10'd43: data = 2'd1;
		10'd44: data = 2'd2;
		10'd45: data = 2'd2;
		10'd46: data = 2'd0;
		10'd47: data = 2'd0;
		10'd48: data = 2'd2;
		10'd49: data = 2'd2;
		10'd50: data = 2'd0;
		10'd51: data = 2'd0;
		10'd52: data = 2'd2;
		10'd53: data = 2'd1;
		10'd54: data = 2'd1;
		10'd55: data = 2'd0;
		10'd56: data = 2'd2;
		10'd57: data = 2'd2;
		10'd58: data = 2'd0;
		10'd59: data = 2'd0;
		10'd60: data = 2'd2;
		10'd61: data = 2'd2;
		10'd62: data = 2'd0;
		10'd63: data = 2'd0;
		10'd64: data = 2'd2;
		10'd65: data = 2'd1;
		10'd66: data = 2'd0;
		10'd67: data = 2'd1;
		10'd68: data = 2'd2;
		10'd69: data = 2'd0;
		10'd70: data = 2'd0;
		10'd71: data = 2'd1;
		10'd72: data = 2'd0;
		10'd73: data = 2'd0;
		10'd74: data = 2'd0;
		10'd75: data = 2'd1;
		10'd76: data = 2'd0;
		10'd77: data = 2'd0;
		10'd78: data = 2'd1;
		10'd79: data = 2'd1;
		10'd80: data = 2'd0;
		10'd81: data = 2'd0;
		10'd82: data = 2'd0;
		10'd83: data = 2'd1;
		10'd84: data = 2'd1;
		10'd85: data = 2'd0;
		10'd86: data = 2'd1;
		10'd87: data = 2'd0;
		10'd88: data = 2'd1;
		10'd89: data = 2'd0;
		10'd90: data = 2'd0;
		10'd91: data = 2'd0;
		10'd92: data = 2'd2;
		10'd93: data = 2'd1;
		10'd94: data = 2'd1;
		10'd95: data = 2'd0;
		10'd96: data = 2'd2;
		10'd97: data = 2'd1;
		10'd98: data = 2'd0;
		10'd99: data = 2'd1;
		10'd100: data = 2'd2;
		10'd101: data = 2'd1;
		10'd102: data = 2'd0;
		10'd103: data = 2'd1;
		10'd104: data = 2'd2;
		10'd105: data = 2'd1;
		10'd106: data = 2'd0;
		10'd107: data = 2'd0;
		10'd108: data = 2'd2;
		10'd109: data = 2'd0;
		10'd110: data = 2'd0;
		10'd111: data = 2'd0;
		10'd112: data = 2'd2;
		10'd113: data = 2'd0;
		10'd114: data = 2'd1;
		10'd115: data = 2'd0;
		10'd116: data = 2'd2;
		10'd117: data = 2'd2;
		10'd118: data = 2'd0;
		10'd119: data = 2'd0;
		10'd120: data = 2'd2;
		10'd121: data = 2'd2;
		10'd122: data = 2'd0;
		10'd123: data = 2'd0;
		10'd124: data = 2'd2;
		10'd125: data = 2'd2;
		10'd126: data = 2'd1;
		10'd127: data = 2'd0;
		10'd128: data = 2'd2;
		10'd129: data = 2'd1;
		10'd130: data = 2'd0;
		10'd131: data = 2'd1;
		10'd132: data = 2'd2;
		10'd133: data = 2'd0;
		10'd134: data = 2'd0;
		10'd135: data = 2'd1;
		10'd136: data = 2'd0;
		10'd137: data = 2'd0;
		10'd138: data = 2'd0;
		10'd139: data = 2'd1;
		10'd140: data = 2'd0;
		10'd141: data = 2'd0;
		10'd142: data = 2'd0;
		10'd143: data = 2'd1;
		10'd144: data = 2'd1;
		10'd145: data = 2'd0;
		10'd146: data = 2'd0;
		10'd147: data = 2'd0;
		10'd148: data = 2'd1;
		10'd149: data = 2'd0;
		10'd150: data = 2'd0;
		10'd151: data = 2'd1;
		10'd152: data = 2'd0;
		10'd153: data = 2'd0;
		10'd154: data = 2'd0;
		10'd155: data = 2'd0;
		10'd156: data = 2'd2;
		10'd157: data = 2'd0;
		10'd158: data = 2'd0;
		10'd159: data = 2'd0;
		10'd160: data = 2'd2;
		10'd161: data = 2'd1;
		10'd162: data = 2'd0;
		10'd163: data = 2'd1;
		10'd164: data = 2'd2;
		10'd165: data = 2'd0;
		10'd166: data = 2'd0;
		10'd167: data = 2'd1;
		10'd168: data = 2'd2;
		10'd169: data = 2'd0;
		10'd170: data = 2'd1;
		10'd171: data = 2'd0;
		10'd172: data = 2'd1;
		10'd173: data = 2'd0;
		10'd174: data = 2'd1;
		10'd175: data = 2'd0;
		10'd176: data = 2'd1;
		10'd177: data = 2'd1;
		10'd178: data = 2'd0;
		10'd179: data = 2'd0;
		10'd180: data = 2'd1;
		10'd181: data = 2'd1;
		10'd182: data = 2'd0;
		10'd183: data = 2'd0;
		10'd184: data = 2'd2;
		10'd185: data = 2'd2;
		10'd186: data = 2'd0;
		10'd187: data = 2'd0;
		10'd188: data = 2'd1;
		10'd189: data = 2'd2;
		10'd190: data = 2'd0;
		10'd191: data = 2'd0;
		10'd192: data = 2'd2;
		10'd193: data = 2'd1;
		10'd194: data = 2'd0;
		10'd195: data = 2'd2;
		10'd196: data = 2'd2;
		10'd197: data = 2'd0;
		10'd198: data = 2'd0;
		10'd199: data = 2'd1;
		10'd200: data = 2'd0;
		10'd201: data = 2'd1;
		10'd202: data = 2'd0;
		10'd203: data = 2'd1;
		10'd204: data = 2'd0;
		10'd205: data = 2'd0;
		10'd206: data = 2'd0;
		10'd207: data = 2'd1;
		10'd208: data = 2'd1;
		10'd209: data = 2'd1;
		10'd210: data = 2'd0;
		10'd211: data = 2'd0;
		10'd212: data = 2'd1;
		10'd213: data = 2'd0;
		10'd214: data = 2'd0;
		10'd215: data = 2'd0;
		10'd216: data = 2'd0;
		10'd217: data = 2'd0;
		10'd218: data = 2'd1;
		10'd219: data = 2'd1;
		10'd220: data = 2'd2;
		10'd221: data = 2'd0;
		10'd222: data = 2'd0;
		10'd223: data = 2'd0;
		10'd224: data = 2'd2;
		10'd225: data = 2'd0;
		10'd226: data = 2'd0;
		10'd227: data = 2'd1;
		10'd228: data = 2'd2;
		10'd229: data = 2'd0;
		10'd230: data = 2'd0;
		10'd231: data = 2'd0;
		10'd232: data = 2'd1;
		10'd233: data = 2'd0;
		10'd234: data = 2'd0;
		10'd235: data = 2'd0;
		10'd236: data = 2'd1;
		10'd237: data = 2'd0;
		10'd238: data = 2'd0;
		10'd239: data = 2'd0;
		10'd240: data = 2'd0;
		10'd241: data = 2'd1;
		10'd242: data = 2'd0;
		10'd243: data = 2'd0;
		10'd244: data = 2'd1;
		10'd245: data = 2'd1;
		10'd246: data = 2'd0;
		10'd247: data = 2'd0;
		10'd248: data = 2'd1;
		10'd249: data = 2'd1;
		10'd250: data = 2'd0;
		10'd251: data = 2'd0;
		10'd252: data = 2'd1;
		10'd253: data = 2'd0;
		10'd254: data = 2'd0;
		10'd255: data = 2'd0;
		10'd256: data = 2'd2;
		10'd257: data = 2'd2;
		10'd258: data = 2'd0;
		10'd259: data = 2'd1;
		10'd260: data = 2'd2;
		10'd261: data = 2'd1;
		10'd262: data = 2'd1;
		10'd263: data = 2'd1;
		10'd264: data = 2'd0;
		10'd265: data = 2'd0;
		10'd266: data = 2'd0;
		10'd267: data = 2'd1;
		10'd268: data = 2'd0;
		10'd269: data = 2'd2;
		10'd270: data = 2'd0;
		10'd271: data = 2'd0;
		10'd272: data = 2'd0;
		10'd273: data = 2'd1;
		10'd274: data = 2'd0;
		10'd275: data = 2'd0;
		10'd276: data = 2'd1;
		10'd277: data = 2'd0;
		10'd278: data = 2'd0;
		10'd279: data = 2'd0;
		10'd280: data = 2'd0;
		10'd281: data = 2'd0;
		10'd282: data = 2'd0;
		10'd283: data = 2'd0;
		10'd284: data = 2'd0;
		10'd285: data = 2'd0;
		10'd286: data = 2'd0;
		10'd287: data = 2'd1;
		10'd288: data = 2'd0;
		10'd289: data = 2'd0;
		10'd290: data = 2'd0;
		10'd291: data = 2'd0;
		10'd292: data = 2'd0;
		10'd293: data = 2'd0;
		10'd294: data = 2'd0;
		10'd295: data = 2'd0;
		10'd296: data = 2'd2;
		10'd297: data = 2'd0;
		10'd298: data = 2'd1;
		10'd299: data = 2'd0;
		10'd300: data = 2'd1;
		10'd301: data = 2'd0;
		10'd302: data = 2'd0;
		10'd303: data = 2'd0;
		10'd304: data = 2'd1;
		10'd305: data = 2'd0;
		10'd306: data = 2'd0;
		10'd307: data = 2'd0;
		10'd308: data = 2'd0;
		10'd309: data = 2'd1;
		10'd310: data = 2'd1;
		10'd311: data = 2'd0;
		10'd312: data = 2'd1;
		10'd313: data = 2'd1;
		10'd314: data = 2'd0;
		10'd315: data = 2'd0;
		10'd316: data = 2'd0;
		10'd317: data = 2'd1;
		10'd318: data = 2'd0;
		10'd319: data = 2'd0;
		10'd320: data = 2'd2;
		10'd321: data = 2'd2;
		10'd322: data = 2'd0;
		10'd323: data = 2'd1;
		10'd324: data = 2'd2;
		10'd325: data = 2'd2;
		10'd326: data = 2'd0;
		10'd327: data = 2'd1;
		10'd328: data = 2'd0;
		10'd329: data = 2'd2;
		10'd330: data = 2'd0;
		10'd331: data = 2'd1;
		10'd332: data = 2'd0;
		10'd333: data = 2'd1;
		10'd334: data = 2'd0;
		10'd335: data = 2'd1;
		10'd336: data = 2'd0;
		10'd337: data = 2'd1;
		10'd338: data = 2'd1;
		10'd339: data = 2'd0;
		10'd340: data = 2'd1;
		10'd341: data = 2'd0;
		10'd342: data = 2'd0;
		10'd343: data = 2'd0;
		10'd344: data = 2'd2;
		10'd345: data = 2'd0;
		10'd346: data = 2'd0;
		10'd347: data = 2'd0;
		10'd348: data = 2'd1;
		10'd349: data = 2'd0;
		10'd350: data = 2'd0;
		10'd351: data = 2'd0;
		10'd352: data = 2'd2;
		10'd353: data = 2'd0;
		10'd354: data = 2'd0;
		10'd355: data = 2'd0;
		10'd356: data = 2'd1;
		10'd357: data = 2'd0;
		10'd358: data = 2'd0;
		10'd359: data = 2'd0;
		10'd360: data = 2'd1;
		10'd361: data = 2'd0;
		10'd362: data = 2'd0;
		10'd363: data = 2'd0;
		10'd364: data = 2'd1;
		10'd365: data = 2'd1;
		10'd366: data = 2'd1;
		10'd367: data = 2'd0;
		10'd368: data = 2'd1;
		10'd369: data = 2'd1;
		10'd370: data = 2'd1;
		10'd371: data = 2'd0;
		10'd372: data = 2'd1;
		10'd373: data = 2'd0;
		10'd374: data = 2'd0;
		10'd375: data = 2'd0;
		10'd376: data = 2'd0;
		10'd377: data = 2'd1;
		10'd378: data = 2'd0;
		10'd379: data = 2'd0;
		10'd380: data = 2'd1;
		10'd381: data = 2'd1;
		10'd382: data = 2'd1;
		10'd383: data = 2'd0;
		10'd384: data = 2'd2;
		10'd385: data = 2'd2;
		10'd386: data = 2'd0;
		10'd387: data = 2'd1;
		10'd388: data = 2'd2;
		10'd389: data = 2'd1;
		10'd390: data = 2'd0;
		10'd391: data = 2'd1;
		10'd392: data = 2'd1;
		10'd393: data = 2'd0;
		10'd394: data = 2'd1;
		10'd395: data = 2'd0;
		10'd396: data = 2'd0;
		10'd397: data = 2'd1;
		10'd398: data = 2'd0;
		10'd399: data = 2'd0;
		10'd400: data = 2'd0;
		10'd401: data = 2'd0;
		10'd402: data = 2'd0;
		10'd403: data = 2'd1;
		10'd404: data = 2'd0;
		10'd405: data = 2'd0;
		10'd406: data = 2'd0;
		10'd407: data = 2'd0;
		10'd408: data = 2'd1;
		10'd409: data = 2'd0;
		10'd410: data = 2'd0;
		10'd411: data = 2'd0;
		10'd412: data = 2'd1;
		10'd413: data = 2'd0;
		10'd414: data = 2'd0;
		10'd415: data = 2'd0;
		10'd416: data = 2'd1;
		10'd417: data = 2'd0;
		10'd418: data = 2'd0;
		10'd419: data = 2'd0;
		10'd420: data = 2'd1;
		10'd421: data = 2'd0;
		10'd422: data = 2'd0;
		10'd423: data = 2'd0;
		10'd424: data = 2'd1;
		10'd425: data = 2'd0;
		10'd426: data = 2'd0;
		10'd427: data = 2'd0;
		10'd428: data = 2'd1;
		10'd429: data = 2'd0;
		10'd430: data = 2'd0;
		10'd431: data = 2'd0;
		10'd432: data = 2'd1;
		10'd433: data = 2'd1;
		10'd434: data = 2'd0;
		10'd435: data = 2'd0;
		10'd436: data = 2'd1;
		10'd437: data = 2'd1;
		10'd438: data = 2'd0;
		10'd439: data = 2'd0;
		10'd440: data = 2'd1;
		10'd441: data = 2'd1;
		10'd442: data = 2'd0;
		10'd443: data = 2'd0;
		10'd444: data = 2'd0;
		10'd445: data = 2'd1;
		10'd446: data = 2'd1;
		10'd447: data = 2'd0;
		10'd448: data = 2'd2;
		10'd449: data = 2'd2;
		10'd450: data = 2'd1;
		10'd451: data = 2'd1;
		10'd452: data = 2'd2;
		10'd453: data = 2'd0;
		10'd454: data = 2'd0;
		10'd455: data = 2'd1;
		10'd456: data = 2'd1;
		10'd457: data = 2'd1;
		10'd458: data = 2'd0;
		10'd459: data = 2'd0;
		10'd460: data = 2'd0;
		10'd461: data = 2'd0;
		10'd462: data = 2'd0;
		10'd463: data = 2'd0;
		10'd464: data = 2'd0;
		10'd465: data = 2'd0;
		10'd466: data = 2'd0;
		10'd467: data = 2'd0;
		10'd468: data = 2'd1;
		10'd469: data = 2'd0;
		10'd470: data = 2'd0;
		10'd471: data = 2'd1;
		10'd472: data = 2'd1;
		10'd473: data = 2'd0;
		10'd474: data = 2'd0;
		10'd475: data = 2'd0;
		10'd476: data = 2'd0;
		10'd477: data = 2'd0;
		10'd478: data = 2'd0;
		10'd479: data = 2'd0;
		10'd480: data = 2'd1;
		10'd481: data = 2'd0;
		10'd482: data = 2'd0;
		10'd483: data = 2'd0;
		10'd484: data = 2'd0;
		10'd485: data = 2'd0;
		10'd486: data = 2'd0;
		10'd487: data = 2'd0;
		10'd488: data = 2'd1;
		10'd489: data = 2'd0;
		10'd490: data = 2'd0;
		10'd491: data = 2'd0;
		10'd492: data = 2'd1;
		10'd493: data = 2'd1;
		10'd494: data = 2'd1;
		10'd495: data = 2'd0;
		10'd496: data = 2'd1;
		10'd497: data = 2'd1;
		10'd498: data = 2'd0;
		10'd499: data = 2'd0;
		10'd500: data = 2'd1;
		10'd501: data = 2'd1;
		10'd502: data = 2'd0;
		10'd503: data = 2'd0;
		10'd504: data = 2'd0;
		10'd505: data = 2'd1;
		10'd506: data = 2'd1;
		10'd507: data = 2'd0;
		10'd508: data = 2'd1;
		10'd509: data = 2'd1;
		10'd510: data = 2'd1;
		10'd511: data = 2'd0;
		10'd512: data = 2'd2;
		10'd513: data = 2'd2;
		10'd514: data = 2'd0;
		10'd515: data = 2'd2;
		10'd516: data = 2'd2;
		10'd517: data = 2'd2;
		10'd518: data = 2'd0;
		10'd519: data = 2'd1;
		10'd520: data = 2'd2;
		10'd521: data = 2'd0;
		10'd522: data = 2'd0;
		10'd523: data = 2'd0;
		10'd524: data = 2'd0;
		10'd525: data = 2'd1;
		10'd526: data = 2'd1;
		10'd527: data = 2'd1;
		10'd528: data = 2'd1;
		10'd529: data = 2'd1;
		10'd530: data = 2'd0;
		10'd531: data = 2'd0;
		10'd532: data = 2'd0;
		10'd533: data = 2'd0;
		10'd534: data = 2'd0;
		10'd535: data = 2'd0;
		10'd536: data = 2'd1;
		10'd537: data = 2'd0;
		10'd538: data = 2'd0;
		10'd539: data = 2'd0;
		10'd540: data = 2'd1;
		10'd541: data = 2'd0;
		10'd542: data = 2'd0;
		10'd543: data = 2'd0;
		10'd544: data = 2'd0;
		10'd545: data = 2'd0;
		10'd546: data = 2'd0;
		10'd547: data = 2'd0;
		10'd548: data = 2'd0;
		10'd549: data = 2'd0;
		10'd550: data = 2'd0;
		10'd551: data = 2'd0;
		10'd552: data = 2'd0;
		10'd553: data = 2'd1;
		10'd554: data = 2'd0;
		10'd555: data = 2'd0;
		10'd556: data = 2'd1;
		10'd557: data = 2'd0;
		10'd558: data = 2'd0;
		10'd559: data = 2'd0;
		10'd560: data = 2'd1;
		10'd561: data = 2'd0;
		10'd562: data = 2'd0;
		10'd563: data = 2'd0;
		10'd564: data = 2'd1;
		10'd565: data = 2'd1;
		10'd566: data = 2'd0;
		10'd567: data = 2'd0;
		10'd568: data = 2'd1;
		10'd569: data = 2'd1;
		10'd570: data = 2'd1;
		10'd571: data = 2'd0;
		10'd572: data = 2'd1;
		10'd573: data = 2'd1;
		10'd574: data = 2'd1;
		10'd575: data = 2'd0;
		10'd576: data = 2'd2;
		10'd577: data = 2'd2;
		10'd578: data = 2'd0;
		10'd579: data = 2'd1;
		10'd580: data = 2'd2;
		10'd581: data = 2'd2;
		10'd582: data = 2'd1;
		10'd583: data = 2'd1;
		10'd584: data = 2'd1;
		10'd585: data = 2'd1;
		10'd586: data = 2'd0;
		10'd587: data = 2'd1;
		10'd588: data = 2'd1;
		10'd589: data = 2'd0;
		10'd590: data = 2'd0;
		10'd591: data = 2'd0;
		10'd592: data = 2'd1;
		10'd593: data = 2'd0;
		10'd594: data = 2'd0;
		10'd595: data = 2'd1;
		10'd596: data = 2'd1;
		10'd597: data = 2'd1;
		10'd598: data = 2'd0;
		10'd599: data = 2'd0;
		10'd600: data = 2'd0;
		10'd601: data = 2'd0;
		10'd602: data = 2'd0;
		10'd603: data = 2'd0;
		10'd604: data = 2'd0;
		10'd605: data = 2'd0;
		10'd606: data = 2'd0;
		10'd607: data = 2'd0;
		10'd608: data = 2'd0;
		10'd609: data = 2'd0;
		10'd610: data = 2'd0;
		10'd611: data = 2'd0;
		10'd612: data = 2'd0;
		10'd613: data = 2'd1;
		10'd614: data = 2'd0;
		10'd615: data = 2'd0;
		10'd616: data = 2'd0;
		10'd617: data = 2'd0;
		10'd618: data = 2'd0;
		10'd619: data = 2'd0;
		10'd620: data = 2'd0;
		10'd621: data = 2'd1;
		10'd622: data = 2'd0;
		10'd623: data = 2'd0;
		10'd624: data = 2'd1;
		10'd625: data = 2'd1;
		10'd626: data = 2'd0;
		10'd627: data = 2'd0;
		10'd628: data = 2'd1;
		10'd629: data = 2'd1;
		10'd630: data = 2'd0;
		10'd631: data = 2'd0;
		10'd632: data = 2'd1;
		10'd633: data = 2'd1;
		10'd634: data = 2'd0;
		10'd635: data = 2'd0;
		10'd636: data = 2'd1;
		10'd637: data = 2'd1;
		10'd638: data = 2'd1;
		10'd639: data = 2'd0;
		10'd640: data = 2'd2;
		10'd641: data = 2'd2;
		10'd642: data = 2'd1;
		10'd643: data = 2'd1;
		10'd644: data = 2'd2;
		10'd645: data = 2'd2;
		10'd646: data = 2'd0;
		10'd647: data = 2'd1;
		10'd648: data = 2'd2;
		10'd649: data = 2'd1;
		10'd650: data = 2'd0;
		10'd651: data = 2'd1;
		10'd652: data = 2'd2;
		10'd653: data = 2'd0;
		10'd654: data = 2'd0;
		10'd655: data = 2'd0;
		10'd656: data = 2'd0;
		10'd657: data = 2'd0;
		10'd658: data = 2'd0;
		10'd659: data = 2'd1;
		10'd660: data = 2'd0;
		10'd661: data = 2'd0;
		10'd662: data = 2'd0;
		10'd663: data = 2'd0;
		10'd664: data = 2'd1;
		10'd665: data = 2'd1;
		10'd666: data = 2'd0;
		10'd667: data = 2'd0;
		10'd668: data = 2'd0;
		10'd669: data = 2'd0;
		10'd670: data = 2'd0;
		10'd671: data = 2'd0;
		10'd672: data = 2'd0;
		10'd673: data = 2'd1;
		10'd674: data = 2'd0;
		10'd675: data = 2'd0;
		10'd676: data = 2'd0;
		10'd677: data = 2'd1;
		10'd678: data = 2'd0;
		10'd679: data = 2'd0;
		10'd680: data = 2'd0;
		10'd681: data = 2'd0;
		10'd682: data = 2'd0;
		10'd683: data = 2'd0;
		10'd684: data = 2'd1;
		10'd685: data = 2'd0;
		10'd686: data = 2'd1;
		10'd687: data = 2'd0;
		10'd688: data = 2'd1;
		10'd689: data = 2'd1;
		10'd690: data = 2'd0;
		10'd691: data = 2'd0;
		10'd692: data = 2'd1;
		10'd693: data = 2'd1;
		10'd694: data = 2'd0;
		10'd695: data = 2'd0;
		10'd696: data = 2'd2;
		10'd697: data = 2'd1;
		10'd698: data = 2'd0;
		10'd699: data = 2'd0;
		10'd700: data = 2'd2;
		10'd701: data = 2'd1;
		10'd702: data = 2'd1;
		10'd703: data = 2'd0;
		10'd704: data = 2'd2;
		10'd705: data = 2'd2;
		10'd706: data = 2'd1;
		10'd707: data = 2'd1;
		10'd708: data = 2'd2;
		10'd709: data = 2'd2;
		10'd710: data = 2'd0;
		10'd711: data = 2'd1;
		10'd712: data = 2'd2;
		10'd713: data = 2'd2;
		10'd714: data = 2'd0;
		10'd715: data = 2'd1;
		10'd716: data = 2'd2;
		10'd717: data = 2'd1;
		10'd718: data = 2'd0;
		10'd719: data = 2'd1;
		10'd720: data = 2'd2;
		10'd721: data = 2'd0;
		10'd722: data = 2'd0;
		10'd723: data = 2'd0;
		10'd724: data = 2'd0;
		10'd725: data = 2'd0;
		10'd726: data = 2'd0;
		10'd727: data = 2'd0;
		10'd728: data = 2'd0;
		10'd729: data = 2'd0;
		10'd730: data = 2'd0;
		10'd731: data = 2'd0;
		10'd732: data = 2'd0;
		10'd733: data = 2'd1;
		10'd734: data = 2'd0;
		10'd735: data = 2'd0;
		10'd736: data = 2'd0;
		10'd737: data = 2'd1;
		10'd738: data = 2'd0;
		10'd739: data = 2'd0;
		10'd740: data = 2'd0;
		10'd741: data = 2'd0;
		10'd742: data = 2'd0;
		10'd743: data = 2'd0;
		10'd744: data = 2'd0;
		10'd745: data = 2'd0;
		10'd746: data = 2'd0;
		10'd747: data = 2'd0;
		10'd748: data = 2'd1;
		10'd749: data = 2'd0;
		10'd750: data = 2'd0;
		10'd751: data = 2'd0;
		10'd752: data = 2'd1;
		10'd753: data = 2'd1;
		10'd754: data = 2'd1;
		10'd755: data = 2'd0;
		10'd756: data = 2'd2;
		10'd757: data = 2'd1;
		10'd758: data = 2'd0;
		10'd759: data = 2'd0;
		10'd760: data = 2'd1;
		10'd761: data = 2'd1;
		10'd762: data = 2'd0;
		10'd763: data = 2'd0;
		10'd764: data = 2'd0;
		10'd765: data = 2'd1;
		10'd766: data = 2'd0;
		10'd767: data = 2'd0;
		10'd768: data = 2'd2;
		10'd769: data = 2'd2;
		10'd770: data = 2'd2;
		10'd771: data = 2'd1;
		10'd772: data = 2'd2;
		10'd773: data = 2'd2;
		10'd774: data = 2'd1;
		10'd775: data = 2'd1;
		10'd776: data = 2'd2;
		10'd777: data = 2'd2;
		10'd778: data = 2'd0;
		10'd779: data = 2'd1;
		10'd780: data = 2'd2;
		10'd781: data = 2'd1;
		10'd782: data = 2'd0;
		10'd783: data = 2'd1;
		10'd784: data = 2'd1;
		10'd785: data = 2'd1;
		10'd786: data = 2'd0;
		10'd787: data = 2'd0;
		10'd788: data = 2'd1;
		10'd789: data = 2'd0;
		10'd790: data = 2'd0;
		10'd791: data = 2'd0;
		10'd792: data = 2'd1;
		10'd793: data = 2'd0;
		10'd794: data = 2'd0;
		10'd795: data = 2'd0;
		10'd796: data = 2'd0;
		10'd797: data = 2'd1;
		10'd798: data = 2'd0;
		10'd799: data = 2'd0;
		10'd800: data = 2'd0;
		10'd801: data = 2'd0;
		10'd802: data = 2'd0;
		10'd803: data = 2'd0;
		10'd804: data = 2'd0;
		10'd805: data = 2'd0;
		10'd806: data = 2'd0;
		10'd807: data = 2'd0;
		10'd808: data = 2'd1;
		10'd809: data = 2'd0;
		10'd810: data = 2'd0;
		10'd811: data = 2'd0;
		10'd812: data = 2'd1;
		10'd813: data = 2'd1;
		10'd814: data = 2'd0;
		10'd815: data = 2'd0;
		10'd816: data = 2'd1;
		10'd817: data = 2'd1;
		10'd818: data = 2'd1;
		10'd819: data = 2'd0;
		10'd820: data = 2'd0;
		10'd821: data = 2'd1;
		10'd822: data = 2'd1;
		10'd823: data = 2'd0;
		10'd824: data = 2'd0;
		10'd825: data = 2'd2;
		10'd826: data = 2'd0;
		10'd827: data = 2'd0;
		10'd828: data = 2'd1;
		10'd829: data = 2'd2;
		10'd830: data = 2'd0;
		10'd831: data = 2'd0;
		10'd832: data = 2'd2;
		10'd833: data = 2'd2;
		10'd834: data = 2'd2;
		10'd835: data = 2'd0;
		10'd836: data = 2'd2;
		10'd837: data = 2'd2;
		10'd838: data = 2'd1;
		10'd839: data = 2'd1;
		10'd840: data = 2'd2;
		10'd841: data = 2'd2;
		10'd842: data = 2'd0;
		10'd843: data = 2'd1;
		10'd844: data = 2'd0;
		10'd845: data = 2'd2;
		10'd846: data = 2'd0;
		10'd847: data = 2'd0;
		10'd848: data = 2'd0;
		10'd849: data = 2'd1;
		10'd850: data = 2'd1;
		10'd851: data = 2'd0;
		10'd852: data = 2'd0;
		10'd853: data = 2'd1;
		10'd854: data = 2'd1;
		10'd855: data = 2'd0;
		10'd856: data = 2'd1;
		10'd857: data = 2'd1;
		10'd858: data = 2'd0;
		10'd859: data = 2'd0;
		10'd860: data = 2'd0;
		10'd861: data = 2'd1;
		10'd862: data = 2'd0;
		10'd863: data = 2'd0;
		10'd864: data = 2'd0;
		10'd865: data = 2'd1;
		10'd866: data = 2'd0;
		10'd867: data = 2'd0;
		10'd868: data = 2'd0;
		10'd869: data = 2'd0;
		10'd870: data = 2'd0;
		10'd871: data = 2'd0;
		10'd872: data = 2'd0;
		10'd873: data = 2'd1;
		10'd874: data = 2'd0;
		10'd875: data = 2'd0;
		10'd876: data = 2'd1;
		10'd877: data = 2'd1;
		10'd878: data = 2'd1;
		10'd879: data = 2'd0;
		10'd880: data = 2'd2;
		10'd881: data = 2'd1;
		10'd882: data = 2'd0;
		10'd883: data = 2'd0;
		10'd884: data = 2'd2;
		10'd885: data = 2'd2;
		10'd886: data = 2'd0;
		10'd887: data = 2'd0;
		10'd888: data = 2'd2;
		10'd889: data = 2'd2;
		10'd890: data = 2'd1;
		10'd891: data = 2'd0;
		10'd892: data = 2'd2;
		10'd893: data = 2'd2;
		10'd894: data = 2'd1;
		10'd895: data = 2'd0;
		10'd896: data = 2'd2;
		10'd897: data = 2'd2;
		10'd898: data = 2'd2;
		10'd899: data = 2'd1;
		10'd900: data = 2'd1;
		10'd901: data = 2'd2;
		10'd902: data = 2'd2;
		10'd903: data = 2'd0;
		10'd904: data = 2'd0;
		10'd905: data = 2'd2;
		10'd906: data = 2'd1;
		10'd907: data = 2'd0;
		10'd908: data = 2'd0;
		10'd909: data = 2'd2;
		10'd910: data = 2'd1;
		10'd911: data = 2'd0;
		10'd912: data = 2'd0;
		10'd913: data = 2'd2;
		10'd914: data = 2'd1;
		10'd915: data = 2'd0;
		10'd916: data = 2'd0;
		10'd917: data = 2'd1;
		10'd918: data = 2'd0;
		10'd919: data = 2'd0;
		10'd920: data = 2'd1;
		10'd921: data = 2'd1;
		10'd922: data = 2'd0;
		10'd923: data = 2'd0;
		10'd924: data = 2'd0;
		10'd925: data = 2'd0;
		10'd926: data = 2'd0;
		10'd927: data = 2'd0;
		10'd928: data = 2'd0;
		10'd929: data = 2'd1;
		10'd930: data = 2'd0;
		10'd931: data = 2'd0;
		10'd932: data = 2'd1;
		10'd933: data = 2'd2;
		10'd934: data = 2'd0;
		10'd935: data = 2'd0;
		10'd936: data = 2'd1;
		10'd937: data = 2'd2;
		10'd938: data = 2'd0;
		10'd939: data = 2'd0;
		10'd940: data = 2'd2;
		10'd941: data = 2'd2;
		10'd942: data = 2'd0;
		10'd943: data = 2'd0;
		10'd944: data = 2'd2;
		10'd945: data = 2'd2;
		10'd946: data = 2'd1;
		10'd947: data = 2'd0;
		10'd948: data = 2'd2;
		10'd949: data = 2'd1;
		10'd950: data = 2'd0;
		10'd951: data = 2'd0;
		10'd952: data = 2'd2;
		10'd953: data = 2'd2;
		10'd954: data = 2'd0;
		10'd955: data = 2'd0;
		10'd956: data = 2'd2;
		10'd957: data = 2'd2;
		10'd958: data = 2'd1;
		10'd959: data = 2'd0;
		10'd960: data = 2'd2;
		10'd961: data = 2'd2;
		10'd962: data = 2'd2;
		10'd963: data = 2'd1;
		10'd964: data = 2'd1;
		10'd965: data = 2'd2;
		10'd966: data = 2'd2;
		10'd967: data = 2'd1;
		10'd968: data = 2'd0;
		10'd969: data = 2'd2;
		10'd970: data = 2'd2;
		10'd971: data = 2'd0;
		10'd972: data = 2'd0;
		10'd973: data = 2'd2;
		10'd974: data = 2'd2;
		10'd975: data = 2'd0;
		10'd976: data = 2'd0;
		10'd977: data = 2'd2;
		10'd978: data = 2'd2;
		10'd979: data = 2'd0;
		10'd980: data = 2'd0;
		10'd981: data = 2'd2;
		10'd982: data = 2'd1;
		10'd983: data = 2'd0;
		10'd984: data = 2'd0;
		10'd985: data = 2'd2;
		10'd986: data = 2'd1;
		10'd987: data = 2'd0;
		10'd988: data = 2'd0;
		10'd989: data = 2'd1;
		10'd990: data = 2'd1;
		10'd991: data = 2'd0;
		10'd992: data = 2'd1;
		10'd993: data = 2'd1;
		10'd994: data = 2'd0;
		10'd995: data = 2'd0;
		10'd996: data = 2'd1;
		10'd997: data = 2'd2;
		10'd998: data = 2'd1;
		10'd999: data = 2'd0;
		10'd1000: data = 2'd1;
		10'd1001: data = 2'd1;
		10'd1002: data = 2'd0;
		10'd1003: data = 2'd0;
		10'd1004: data = 2'd2;
		10'd1005: data = 2'd1;
		10'd1006: data = 2'd0;
		10'd1007: data = 2'd0;
		10'd1008: data = 2'd2;
		10'd1009: data = 2'd1;
		10'd1010: data = 2'd1;
		10'd1011: data = 2'd0;
		10'd1012: data = 2'd2;
		10'd1013: data = 2'd2;
		10'd1014: data = 2'd1;
		10'd1015: data = 2'd0;
		10'd1016: data = 2'd2;
		10'd1017: data = 2'd2;
		10'd1018: data = 2'd2;
		10'd1019: data = 2'd0;
		10'd1020: data = 2'd0;
		10'd1021: data = 2'd2;
		10'd1022: data = 2'd2;
		10'd1023: data = 2'd0;
		default: data = 2'd0;
	endcase
end
endmodule

module layer1_N4(address, data);
input wire [11:0] address;
output reg [3:0] data;

wire [5:0] i; layer1_N4_idx_1 idx_1_inst(address[11:2], i);
wire [1:0] t; layer1_N4_rsh_1 rsh_1_inst(address[11:2], t);
wire [3:0] b; layer1_N4_2 layer1_N4_2_inst(address[11:2], b);
wire [2:0] u; layer1_N4_ust_1 ust_1_inst({i, address[1:0]}, u);

always @(*) begin
	data = (u >> t) + b;
end
endmodule
